magic
tech sky130A
magscale 1 2
timestamp 1657014066
<< viali >>
rect 77125 37417 77159 37451
rect 77861 37417 77895 37451
rect 20361 37281 20395 37315
rect 22201 37281 22235 37315
rect 24685 37281 24719 37315
rect 26065 37281 26099 37315
rect 27997 37281 28031 37315
rect 29561 37281 29595 37315
rect 32137 37281 32171 37315
rect 35265 37281 35299 37315
rect 37289 37281 37323 37315
rect 39865 37281 39899 37315
rect 42901 37281 42935 37315
rect 45017 37281 45051 37315
rect 1409 37213 1443 37247
rect 2881 37213 2915 37247
rect 4813 37213 4847 37247
rect 6745 37213 6779 37247
rect 8953 37213 8987 37247
rect 10517 37213 10551 37247
rect 12449 37213 12483 37247
rect 14381 37213 14415 37247
rect 16681 37213 16715 37247
rect 18153 37213 18187 37247
rect 20177 37213 20211 37247
rect 22017 37213 22051 37247
rect 24501 37213 24535 37247
rect 25881 37213 25915 37247
rect 27813 37213 27847 37247
rect 29837 37213 29871 37247
rect 32413 37213 32447 37247
rect 35541 37213 35575 37247
rect 37565 37213 37599 37247
rect 40141 37213 40175 37247
rect 43177 37213 43211 37247
rect 45293 37213 45327 37247
rect 46949 37213 46983 37247
rect 48789 37213 48823 37247
rect 50721 37213 50755 37247
rect 52929 37213 52963 37247
rect 54585 37213 54619 37247
rect 56425 37213 56459 37247
rect 58357 37213 58391 37247
rect 60657 37213 60691 37247
rect 62129 37213 62163 37247
rect 64061 37213 64095 37247
rect 65993 37213 66027 37247
rect 68385 37213 68419 37247
rect 69765 37213 69799 37247
rect 71697 37213 71731 37247
rect 73629 37213 73663 37247
rect 75377 37213 75411 37247
rect 76113 37213 76147 37247
rect 76941 37213 76975 37247
rect 77677 37213 77711 37247
rect 1593 37077 1627 37111
rect 3065 37077 3099 37111
rect 4997 37077 5031 37111
rect 6929 37077 6963 37111
rect 9137 37077 9171 37111
rect 10701 37077 10735 37111
rect 12633 37077 12667 37111
rect 14565 37077 14599 37111
rect 16865 37077 16899 37111
rect 18337 37077 18371 37111
rect 46765 37077 46799 37111
rect 48605 37077 48639 37111
rect 50537 37077 50571 37111
rect 52745 37077 52779 37111
rect 54401 37077 54435 37111
rect 56241 37077 56275 37111
rect 58173 37077 58207 37111
rect 60473 37077 60507 37111
rect 61945 37077 61979 37111
rect 63877 37077 63911 37111
rect 65809 37077 65843 37111
rect 68201 37077 68235 37111
rect 69581 37077 69615 37111
rect 71513 37077 71547 37111
rect 73445 37077 73479 37111
rect 75193 37077 75227 37111
rect 75929 37077 75963 37111
rect 73721 36873 73755 36907
rect 74733 36873 74767 36907
rect 75101 36873 75135 36907
rect 77125 36873 77159 36907
rect 33425 36737 33459 36771
rect 41061 36737 41095 36771
rect 76941 36737 76975 36771
rect 77677 36737 77711 36771
rect 33701 36669 33735 36703
rect 41337 36669 41371 36703
rect 73813 36669 73847 36703
rect 73997 36669 74031 36703
rect 75193 36669 75227 36703
rect 75285 36669 75319 36703
rect 77861 36601 77895 36635
rect 73353 36533 73387 36567
rect 73629 36261 73663 36295
rect 73813 36125 73847 36159
rect 77401 36125 77435 36159
rect 77861 36125 77895 36159
rect 77217 35989 77251 36023
rect 78045 35989 78079 36023
rect 71513 35785 71547 35819
rect 72341 35785 72375 35819
rect 72525 35649 72559 35683
rect 77953 35649 77987 35683
rect 71605 35581 71639 35615
rect 71697 35581 71731 35615
rect 71145 35513 71179 35547
rect 77769 35445 77803 35479
rect 77861 35037 77895 35071
rect 78045 34901 78079 34935
rect 69213 34697 69247 34731
rect 69581 34697 69615 34731
rect 70409 34697 70443 34731
rect 77033 34697 77067 34731
rect 69673 34561 69707 34595
rect 70593 34561 70627 34595
rect 77217 34561 77251 34595
rect 77677 34561 77711 34595
rect 69765 34493 69799 34527
rect 77861 34357 77895 34391
rect 76205 34153 76239 34187
rect 76849 34153 76883 34187
rect 68385 34017 68419 34051
rect 77401 34017 77435 34051
rect 68109 33949 68143 33983
rect 76389 33949 76423 33983
rect 77309 33881 77343 33915
rect 67741 33813 67775 33847
rect 68201 33813 68235 33847
rect 77217 33813 77251 33847
rect 72157 33609 72191 33643
rect 77217 33609 77251 33643
rect 77585 33609 77619 33643
rect 68477 33473 68511 33507
rect 71973 33473 72007 33507
rect 77677 33473 77711 33507
rect 77769 33405 77803 33439
rect 68293 33337 68327 33371
rect 78045 32997 78079 33031
rect 77861 32861 77895 32895
rect 65993 32385 66027 32419
rect 77677 32385 77711 32419
rect 65809 32181 65843 32215
rect 77861 32181 77895 32215
rect 65625 31977 65659 32011
rect 66177 31841 66211 31875
rect 62865 31773 62899 31807
rect 63049 31773 63083 31807
rect 64061 31773 64095 31807
rect 64337 31773 64371 31807
rect 65993 31705 66027 31739
rect 66085 31637 66119 31671
rect 61945 31433 61979 31467
rect 63509 31433 63543 31467
rect 63877 31433 63911 31467
rect 63969 31297 64003 31331
rect 77677 31297 77711 31331
rect 62037 31229 62071 31263
rect 62129 31229 62163 31263
rect 64061 31229 64095 31263
rect 61577 31093 61611 31127
rect 77861 31093 77895 31127
rect 62129 30753 62163 30787
rect 62405 30685 62439 30719
rect 58449 30277 58483 30311
rect 77677 30209 77711 30243
rect 58541 30141 58575 30175
rect 58725 30141 58759 30175
rect 60289 30141 60323 30175
rect 60565 30141 60599 30175
rect 77861 30073 77895 30107
rect 58081 30005 58115 30039
rect 60473 29801 60507 29835
rect 58725 29665 58759 29699
rect 61025 29665 61059 29699
rect 59001 29597 59035 29631
rect 77861 29597 77895 29631
rect 60841 29529 60875 29563
rect 60933 29461 60967 29495
rect 78045 29461 78079 29495
rect 77861 28509 77895 28543
rect 78045 28373 78079 28407
rect 56333 28033 56367 28067
rect 56425 27829 56459 27863
rect 55689 27625 55723 27659
rect 54585 27489 54619 27523
rect 56241 27489 56275 27523
rect 54401 27421 54435 27455
rect 56057 27421 56091 27455
rect 77861 27421 77895 27455
rect 54033 27285 54067 27319
rect 54493 27285 54527 27319
rect 56149 27285 56183 27319
rect 78045 27285 78079 27319
rect 54677 27013 54711 27047
rect 77677 26945 77711 26979
rect 54769 26741 54803 26775
rect 77861 26741 77895 26775
rect 52101 26469 52135 26503
rect 52653 26401 52687 26435
rect 52469 26333 52503 26367
rect 53389 26333 53423 26367
rect 52561 26265 52595 26299
rect 53573 26265 53607 26299
rect 77677 25857 77711 25891
rect 77861 25653 77895 25687
rect 50721 25313 50755 25347
rect 50537 25245 50571 25279
rect 51457 25177 51491 25211
rect 50169 25109 50203 25143
rect 50629 25109 50663 25143
rect 51549 25109 51583 25143
rect 48881 24905 48915 24939
rect 48973 24769 49007 24803
rect 77677 24769 77711 24803
rect 49065 24701 49099 24735
rect 48513 24565 48547 24599
rect 77861 24565 77895 24599
rect 49249 24157 49283 24191
rect 49341 24021 49375 24055
rect 49709 23817 49743 23851
rect 49617 23681 49651 23715
rect 77309 23681 77343 23715
rect 77677 23681 77711 23715
rect 77861 23545 77895 23579
rect 47041 23205 47075 23239
rect 77861 23069 77895 23103
rect 46857 23001 46891 23035
rect 77493 22933 77527 22967
rect 78045 22933 78079 22967
rect 44833 22729 44867 22763
rect 46213 22729 46247 22763
rect 46581 22729 46615 22763
rect 44925 22593 44959 22627
rect 49985 22593 50019 22627
rect 45017 22525 45051 22559
rect 46673 22525 46707 22559
rect 46765 22525 46799 22559
rect 44465 22389 44499 22423
rect 50077 22389 50111 22423
rect 45201 22185 45235 22219
rect 40417 22049 40451 22083
rect 43085 22049 43119 22083
rect 40233 21981 40267 22015
rect 42901 21981 42935 22015
rect 43729 21981 43763 22015
rect 45017 21981 45051 22015
rect 77861 21981 77895 22015
rect 42533 21845 42567 21879
rect 42993 21845 43027 21879
rect 43913 21845 43947 21879
rect 78045 21845 78079 21879
rect 40509 20961 40543 20995
rect 41705 20961 41739 20995
rect 40233 20893 40267 20927
rect 41429 20893 41463 20927
rect 77861 20893 77895 20927
rect 77493 20825 77527 20859
rect 39865 20757 39899 20791
rect 40325 20757 40359 20791
rect 41061 20757 41095 20791
rect 41521 20757 41555 20791
rect 78045 20757 78079 20791
rect 41429 20553 41463 20587
rect 39681 20417 39715 20451
rect 41245 20417 41279 20451
rect 50353 20417 50387 20451
rect 77677 20417 77711 20451
rect 50997 20349 51031 20383
rect 39865 20281 39899 20315
rect 77861 20213 77895 20247
rect 77677 19329 77711 19363
rect 77309 19125 77343 19159
rect 77861 19125 77895 19159
rect 37197 18717 37231 18751
rect 37381 18581 37415 18615
rect 37289 18377 37323 18411
rect 37657 18377 37691 18411
rect 77309 18241 77343 18275
rect 77677 18241 77711 18275
rect 37749 18173 37783 18207
rect 37841 18173 37875 18207
rect 77861 18037 77895 18071
rect 36277 17833 36311 17867
rect 34897 17765 34931 17799
rect 35449 17697 35483 17731
rect 36093 17629 36127 17663
rect 77861 17629 77895 17663
rect 35265 17561 35299 17595
rect 35357 17493 35391 17527
rect 78045 17493 78079 17527
rect 33425 17289 33459 17323
rect 36553 17221 36587 17255
rect 36737 17221 36771 17255
rect 34253 17153 34287 17187
rect 33517 17085 33551 17119
rect 33701 17085 33735 17119
rect 33057 17017 33091 17051
rect 34437 17017 34471 17051
rect 31585 16609 31619 16643
rect 31677 16609 31711 16643
rect 31493 16541 31527 16575
rect 77861 16541 77895 16575
rect 31125 16405 31159 16439
rect 78045 16405 78079 16439
rect 29929 16201 29963 16235
rect 32229 16133 32263 16167
rect 30021 15997 30055 16031
rect 30205 15997 30239 16031
rect 29561 15861 29595 15895
rect 32505 15861 32539 15895
rect 14381 15657 14415 15691
rect 30297 15453 30331 15487
rect 77861 15453 77895 15487
rect 14289 15385 14323 15419
rect 30573 15317 30607 15351
rect 78045 15317 78079 15351
rect 14657 15113 14691 15147
rect 16865 15113 16899 15147
rect 18429 15113 18463 15147
rect 13461 14977 13495 15011
rect 15209 14977 15243 15011
rect 16773 14977 16807 15011
rect 18337 14977 18371 15011
rect 14197 14909 14231 14943
rect 15393 14909 15427 14943
rect 14565 14841 14599 14875
rect 13645 14773 13679 14807
rect 14657 14569 14691 14603
rect 16313 14569 16347 14603
rect 14473 14501 14507 14535
rect 16221 14501 16255 14535
rect 17601 14501 17635 14535
rect 18337 14365 18371 14399
rect 27077 14365 27111 14399
rect 77861 14365 77895 14399
rect 14197 14297 14231 14331
rect 15853 14297 15887 14331
rect 17233 14297 17267 14331
rect 27813 14297 27847 14331
rect 17693 14229 17727 14263
rect 18153 14229 18187 14263
rect 27169 14229 27203 14263
rect 28089 14229 28123 14263
rect 78045 14229 78079 14263
rect 14657 14025 14691 14059
rect 27169 14025 27203 14059
rect 27537 14025 27571 14059
rect 14197 13957 14231 13991
rect 77309 13957 77343 13991
rect 77677 13889 77711 13923
rect 27629 13821 27663 13855
rect 27721 13821 27755 13855
rect 14473 13753 14507 13787
rect 77861 13685 77895 13719
rect 26985 13481 27019 13515
rect 25973 13345 26007 13379
rect 25789 13277 25823 13311
rect 26709 13209 26743 13243
rect 25421 13141 25455 13175
rect 25881 13141 25915 13175
rect 77677 12801 77711 12835
rect 77309 12597 77343 12631
rect 77861 12597 77895 12631
rect 24777 12393 24811 12427
rect 23673 12257 23707 12291
rect 23489 12189 23523 12223
rect 24501 12121 24535 12155
rect 23121 12053 23155 12087
rect 23581 12053 23615 12087
rect 20361 11849 20395 11883
rect 21833 11849 21867 11883
rect 22201 11849 22235 11883
rect 23857 11781 23891 11815
rect 77677 11713 77711 11747
rect 20453 11645 20487 11679
rect 20637 11645 20671 11679
rect 22293 11645 22327 11679
rect 22385 11645 22419 11679
rect 77861 11577 77895 11611
rect 19993 11509 20027 11543
rect 24133 11509 24167 11543
rect 78045 11237 78079 11271
rect 23397 11101 23431 11135
rect 23765 11101 23799 11135
rect 77861 11101 77895 11135
rect 77953 10081 77987 10115
rect 77677 10013 77711 10047
rect 8309 9129 8343 9163
rect 9137 9061 9171 9095
rect 8953 8925 8987 8959
rect 77677 8925 77711 8959
rect 8217 8857 8251 8891
rect 77953 8857 77987 8891
rect 8217 8585 8251 8619
rect 10609 8585 10643 8619
rect 8125 8449 8159 8483
rect 9781 8449 9815 8483
rect 10517 8449 10551 8483
rect 8769 8381 8803 8415
rect 9229 8381 9263 8415
rect 9045 8313 9079 8347
rect 9965 8313 9999 8347
rect 8401 8041 8435 8075
rect 9413 8041 9447 8075
rect 10333 8041 10367 8075
rect 8217 7973 8251 8007
rect 9321 7973 9355 8007
rect 10241 7973 10275 8007
rect 77677 7837 77711 7871
rect 7941 7769 7975 7803
rect 8953 7769 8987 7803
rect 9873 7769 9907 7803
rect 77953 7769 77987 7803
rect 9229 7497 9263 7531
rect 9689 7497 9723 7531
rect 8769 7429 8803 7463
rect 9873 7361 9907 7395
rect 77493 7361 77527 7395
rect 77769 7293 77803 7327
rect 9137 7225 9171 7259
rect 77493 6273 77527 6307
rect 77677 6205 77711 6239
rect 77493 5185 77527 5219
rect 77677 5117 77711 5151
rect 77677 4573 77711 4607
rect 77953 4505 77987 4539
rect 77769 4165 77803 4199
rect 77953 4097 77987 4131
rect 9597 3689 9631 3723
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 14473 3485 14507 3519
rect 15853 3485 15887 3519
rect 16497 3485 16531 3519
rect 77677 3485 77711 3519
rect 77953 3417 77987 3451
rect 8217 3349 8251 3383
rect 9781 3349 9815 3383
rect 14289 3349 14323 3383
rect 15669 3349 15703 3383
rect 16313 3349 16347 3383
rect 14013 3145 14047 3179
rect 14381 3145 14415 3179
rect 16221 3145 16255 3179
rect 16681 3145 16715 3179
rect 76941 3145 76975 3179
rect 9321 3077 9355 3111
rect 8401 3009 8435 3043
rect 9137 3009 9171 3043
rect 9597 3009 9631 3043
rect 10057 3009 10091 3043
rect 10241 3009 10275 3043
rect 10701 3009 10735 3043
rect 13737 3009 13771 3043
rect 14565 3009 14599 3043
rect 14749 3009 14783 3043
rect 15301 3009 15335 3043
rect 15393 3009 15427 3043
rect 16865 3009 16899 3043
rect 17693 3009 17727 3043
rect 17877 3009 17911 3043
rect 18521 3009 18555 3043
rect 41337 3009 41371 3043
rect 76849 3009 76883 3043
rect 77493 3009 77527 3043
rect 77769 3009 77803 3043
rect 8953 2941 8987 2975
rect 9413 2941 9447 2975
rect 9873 2941 9907 2975
rect 17049 2941 17083 2975
rect 17509 2941 17543 2975
rect 41061 2941 41095 2975
rect 10517 2873 10551 2907
rect 13553 2873 13587 2907
rect 18245 2873 18279 2907
rect 8217 2805 8251 2839
rect 9781 2805 9815 2839
rect 15577 2805 15611 2839
rect 18337 2805 18371 2839
rect 13369 2601 13403 2635
rect 14289 2601 14323 2635
rect 20085 2601 20119 2635
rect 21925 2601 21959 2635
rect 24409 2601 24443 2635
rect 25789 2601 25823 2635
rect 27721 2601 27755 2635
rect 29561 2601 29595 2635
rect 32137 2601 32171 2635
rect 47823 2601 47857 2635
rect 49065 2601 49099 2635
rect 50721 2601 50755 2635
rect 52929 2601 52963 2635
rect 54585 2601 54619 2635
rect 56425 2601 56459 2635
rect 58357 2601 58391 2635
rect 62129 2601 62163 2635
rect 64061 2601 64095 2635
rect 65993 2601 66027 2635
rect 68385 2601 68419 2635
rect 69765 2601 69799 2635
rect 71697 2601 71731 2635
rect 73629 2601 73663 2635
rect 75285 2601 75319 2635
rect 7481 2533 7515 2567
rect 9505 2465 9539 2499
rect 10149 2465 10183 2499
rect 14657 2465 14691 2499
rect 76757 2465 76791 2499
rect 1409 2397 1443 2431
rect 2881 2397 2915 2431
rect 4813 2397 4847 2431
rect 6745 2397 6779 2431
rect 7665 2397 7699 2431
rect 8125 2397 8159 2431
rect 9873 2397 9907 2431
rect 9965 2397 9999 2431
rect 10609 2397 10643 2431
rect 11713 2397 11747 2431
rect 12449 2397 12483 2431
rect 13553 2397 13587 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 15117 2397 15151 2431
rect 16681 2397 16715 2431
rect 18153 2397 18187 2431
rect 20269 2397 20303 2431
rect 22109 2397 22143 2431
rect 24593 2397 24627 2431
rect 25973 2397 26007 2431
rect 27905 2397 27939 2431
rect 29745 2397 29779 2431
rect 32321 2397 32355 2431
rect 33333 2397 33367 2431
rect 33609 2397 33643 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37289 2397 37323 2431
rect 37565 2397 37599 2431
rect 39865 2397 39899 2431
rect 40141 2397 40175 2431
rect 42901 2397 42935 2431
rect 43177 2397 43211 2431
rect 45017 2397 45051 2431
rect 45293 2397 45327 2431
rect 47593 2397 47627 2431
rect 60749 2397 60783 2431
rect 73445 2397 73479 2431
rect 75101 2397 75135 2431
rect 76573 2397 76607 2431
rect 77493 2397 77527 2431
rect 48973 2329 49007 2363
rect 50629 2329 50663 2363
rect 52837 2329 52871 2363
rect 54493 2329 54527 2363
rect 56333 2329 56367 2363
rect 58265 2329 58299 2363
rect 60565 2329 60599 2363
rect 62037 2329 62071 2363
rect 63969 2329 64003 2363
rect 65901 2329 65935 2363
rect 68293 2329 68327 2363
rect 69673 2329 69707 2363
rect 71605 2329 71639 2363
rect 77769 2329 77803 2363
rect 1593 2261 1627 2295
rect 3065 2261 3099 2295
rect 4997 2261 5031 2295
rect 6929 2261 6963 2295
rect 8309 2261 8343 2295
rect 10793 2261 10827 2295
rect 11529 2261 11563 2295
rect 12633 2261 12667 2295
rect 15301 2261 15335 2295
rect 16865 2261 16899 2295
rect 18337 2261 18371 2295
<< metal1 >>
rect 1104 37562 78844 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 78844 37562
rect 1104 37488 78844 37510
rect 77113 37451 77171 37457
rect 77113 37417 77125 37451
rect 77159 37448 77171 37451
rect 77202 37448 77208 37460
rect 77159 37420 77208 37448
rect 77159 37417 77171 37420
rect 77113 37411 77171 37417
rect 77202 37408 77208 37420
rect 77260 37408 77266 37460
rect 77846 37448 77852 37460
rect 77807 37420 77852 37448
rect 77846 37408 77852 37420
rect 77904 37408 77910 37460
rect 20346 37312 20352 37324
rect 20307 37284 20352 37312
rect 20346 37272 20352 37284
rect 20404 37272 20410 37324
rect 22186 37312 22192 37324
rect 22147 37284 22192 37312
rect 22186 37272 22192 37284
rect 22244 37272 22250 37324
rect 23474 37272 23480 37324
rect 23532 37312 23538 37324
rect 24673 37315 24731 37321
rect 24673 37312 24685 37315
rect 23532 37284 24685 37312
rect 23532 37272 23538 37284
rect 24673 37281 24685 37284
rect 24719 37281 24731 37315
rect 24673 37275 24731 37281
rect 25774 37272 25780 37324
rect 25832 37312 25838 37324
rect 26053 37315 26111 37321
rect 26053 37312 26065 37315
rect 25832 37284 26065 37312
rect 25832 37272 25838 37284
rect 26053 37281 26065 37284
rect 26099 37281 26111 37315
rect 26053 37275 26111 37281
rect 27522 37272 27528 37324
rect 27580 37312 27586 37324
rect 27985 37315 28043 37321
rect 27985 37312 27997 37315
rect 27580 37284 27997 37312
rect 27580 37272 27586 37284
rect 27985 37281 27997 37284
rect 28031 37281 28043 37315
rect 27985 37275 28043 37281
rect 29454 37272 29460 37324
rect 29512 37312 29518 37324
rect 29549 37315 29607 37321
rect 29549 37312 29561 37315
rect 29512 37284 29561 37312
rect 29512 37272 29518 37284
rect 29549 37281 29561 37284
rect 29595 37281 29607 37315
rect 29549 37275 29607 37281
rect 31386 37272 31392 37324
rect 31444 37312 31450 37324
rect 32125 37315 32183 37321
rect 32125 37312 32137 37315
rect 31444 37284 32137 37312
rect 31444 37272 31450 37284
rect 32125 37281 32137 37284
rect 32171 37281 32183 37315
rect 32125 37275 32183 37281
rect 35253 37315 35311 37321
rect 35253 37281 35265 37315
rect 35299 37312 35311 37315
rect 35342 37312 35348 37324
rect 35299 37284 35348 37312
rect 35299 37281 35311 37284
rect 35253 37275 35311 37281
rect 35342 37272 35348 37284
rect 35400 37272 35406 37324
rect 37090 37272 37096 37324
rect 37148 37312 37154 37324
rect 37277 37315 37335 37321
rect 37277 37312 37289 37315
rect 37148 37284 37289 37312
rect 37148 37272 37154 37284
rect 37277 37281 37289 37284
rect 37323 37281 37335 37315
rect 37277 37275 37335 37281
rect 39022 37272 39028 37324
rect 39080 37312 39086 37324
rect 39853 37315 39911 37321
rect 39853 37312 39865 37315
rect 39080 37284 39865 37312
rect 39080 37272 39086 37284
rect 39853 37281 39865 37284
rect 39899 37281 39911 37315
rect 39853 37275 39911 37281
rect 42794 37272 42800 37324
rect 42852 37312 42858 37324
rect 42889 37315 42947 37321
rect 42889 37312 42901 37315
rect 42852 37284 42901 37312
rect 42852 37272 42858 37284
rect 42889 37281 42901 37284
rect 42935 37281 42947 37315
rect 42889 37275 42947 37281
rect 44726 37272 44732 37324
rect 44784 37312 44790 37324
rect 45005 37315 45063 37321
rect 45005 37312 45017 37315
rect 44784 37284 45017 37312
rect 44784 37272 44790 37284
rect 45005 37281 45017 37284
rect 45051 37281 45063 37315
rect 45005 37275 45063 37281
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 2866 37244 2872 37256
rect 2827 37216 2872 37244
rect 2866 37204 2872 37216
rect 2924 37204 2930 37256
rect 4798 37244 4804 37256
rect 4759 37216 4804 37244
rect 4798 37204 4804 37216
rect 4856 37204 4862 37256
rect 6730 37244 6736 37256
rect 6691 37216 6736 37244
rect 6730 37204 6736 37216
rect 6788 37204 6794 37256
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 8941 37247 8999 37253
rect 8941 37244 8953 37247
rect 8352 37216 8953 37244
rect 8352 37204 8358 37216
rect 8941 37213 8953 37216
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 10505 37247 10563 37253
rect 10505 37213 10517 37247
rect 10551 37244 10563 37247
rect 10594 37244 10600 37256
rect 10551 37216 10600 37244
rect 10551 37213 10563 37216
rect 10505 37207 10563 37213
rect 10594 37204 10600 37216
rect 10652 37204 10658 37256
rect 12434 37244 12440 37256
rect 12395 37216 12440 37244
rect 12434 37204 12440 37216
rect 12492 37204 12498 37256
rect 14366 37244 14372 37256
rect 14327 37216 14372 37244
rect 14366 37204 14372 37216
rect 14424 37204 14430 37256
rect 16669 37247 16727 37253
rect 16669 37213 16681 37247
rect 16715 37244 16727 37247
rect 16758 37244 16764 37256
rect 16715 37216 16764 37244
rect 16715 37213 16727 37216
rect 16669 37207 16727 37213
rect 16758 37204 16764 37216
rect 16816 37204 16822 37256
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37244 18199 37247
rect 18414 37244 18420 37256
rect 18187 37216 18420 37244
rect 18187 37213 18199 37216
rect 18141 37207 18199 37213
rect 18414 37204 18420 37216
rect 18472 37204 18478 37256
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 20036 37216 20177 37244
rect 20036 37204 20042 37216
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 20165 37207 20223 37213
rect 21818 37204 21824 37256
rect 21876 37244 21882 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21876 37216 22017 37244
rect 21876 37204 21882 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 23750 37204 23756 37256
rect 23808 37244 23814 37256
rect 24489 37247 24547 37253
rect 24489 37244 24501 37247
rect 23808 37216 24501 37244
rect 23808 37204 23814 37216
rect 24489 37213 24501 37216
rect 24535 37213 24547 37247
rect 24489 37207 24547 37213
rect 25682 37204 25688 37256
rect 25740 37244 25746 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25740 37216 25881 37244
rect 25740 37204 25746 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 27614 37204 27620 37256
rect 27672 37244 27678 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27672 37216 27813 37244
rect 27672 37204 27678 37216
rect 27801 37213 27813 37216
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 29825 37247 29883 37253
rect 29825 37213 29837 37247
rect 29871 37244 29883 37247
rect 29914 37244 29920 37256
rect 29871 37216 29920 37244
rect 29871 37213 29883 37216
rect 29825 37207 29883 37213
rect 29914 37204 29920 37216
rect 29972 37204 29978 37256
rect 32398 37244 32404 37256
rect 32359 37216 32404 37244
rect 32398 37204 32404 37216
rect 32456 37204 32462 37256
rect 35434 37204 35440 37256
rect 35492 37244 35498 37256
rect 35529 37247 35587 37253
rect 35529 37244 35541 37247
rect 35492 37216 35541 37244
rect 35492 37204 35498 37216
rect 35529 37213 35541 37216
rect 35575 37213 35587 37247
rect 35529 37207 35587 37213
rect 37553 37247 37611 37253
rect 37553 37213 37565 37247
rect 37599 37244 37611 37247
rect 37642 37244 37648 37256
rect 37599 37216 37648 37244
rect 37599 37213 37611 37216
rect 37553 37207 37611 37213
rect 37642 37204 37648 37216
rect 37700 37204 37706 37256
rect 40129 37247 40187 37253
rect 40129 37213 40141 37247
rect 40175 37244 40187 37247
rect 40218 37244 40224 37256
rect 40175 37216 40224 37244
rect 40175 37213 40187 37216
rect 40129 37207 40187 37213
rect 40218 37204 40224 37216
rect 40276 37204 40282 37256
rect 43165 37247 43223 37253
rect 43165 37244 43177 37247
rect 42812 37216 43177 37244
rect 42812 37188 42840 37216
rect 43165 37213 43177 37216
rect 43211 37213 43223 37247
rect 43165 37207 43223 37213
rect 44818 37204 44824 37256
rect 44876 37244 44882 37256
rect 45281 37247 45339 37253
rect 45281 37244 45293 37247
rect 44876 37216 45293 37244
rect 44876 37204 44882 37216
rect 45281 37213 45293 37216
rect 45327 37213 45339 37247
rect 45281 37207 45339 37213
rect 46658 37204 46664 37256
rect 46716 37244 46722 37256
rect 46937 37247 46995 37253
rect 46937 37244 46949 37247
rect 46716 37216 46949 37244
rect 46716 37204 46722 37216
rect 46937 37213 46949 37216
rect 46983 37213 46995 37247
rect 46937 37207 46995 37213
rect 48498 37204 48504 37256
rect 48556 37244 48562 37256
rect 48777 37247 48835 37253
rect 48777 37244 48789 37247
rect 48556 37216 48789 37244
rect 48556 37204 48562 37216
rect 48777 37213 48789 37216
rect 48823 37213 48835 37247
rect 48777 37207 48835 37213
rect 50430 37204 50436 37256
rect 50488 37244 50494 37256
rect 50709 37247 50767 37253
rect 50709 37244 50721 37247
rect 50488 37216 50721 37244
rect 50488 37204 50494 37216
rect 50709 37213 50721 37216
rect 50755 37213 50767 37247
rect 50709 37207 50767 37213
rect 52454 37204 52460 37256
rect 52512 37244 52518 37256
rect 52917 37247 52975 37253
rect 52917 37244 52929 37247
rect 52512 37216 52929 37244
rect 52512 37204 52518 37216
rect 52917 37213 52929 37216
rect 52963 37213 52975 37247
rect 52917 37207 52975 37213
rect 54294 37204 54300 37256
rect 54352 37244 54358 37256
rect 54573 37247 54631 37253
rect 54573 37244 54585 37247
rect 54352 37216 54585 37244
rect 54352 37204 54358 37216
rect 54573 37213 54585 37216
rect 54619 37213 54631 37247
rect 54573 37207 54631 37213
rect 56134 37204 56140 37256
rect 56192 37244 56198 37256
rect 56413 37247 56471 37253
rect 56413 37244 56425 37247
rect 56192 37216 56425 37244
rect 56192 37204 56198 37216
rect 56413 37213 56425 37216
rect 56459 37213 56471 37247
rect 56413 37207 56471 37213
rect 58066 37204 58072 37256
rect 58124 37244 58130 37256
rect 58345 37247 58403 37253
rect 58345 37244 58357 37247
rect 58124 37216 58357 37244
rect 58124 37204 58130 37216
rect 58345 37213 58357 37216
rect 58391 37213 58403 37247
rect 58345 37207 58403 37213
rect 59998 37204 60004 37256
rect 60056 37244 60062 37256
rect 60645 37247 60703 37253
rect 60645 37244 60657 37247
rect 60056 37216 60657 37244
rect 60056 37204 60062 37216
rect 60645 37213 60657 37216
rect 60691 37213 60703 37247
rect 60645 37207 60703 37213
rect 61838 37204 61844 37256
rect 61896 37244 61902 37256
rect 62117 37247 62175 37253
rect 62117 37244 62129 37247
rect 61896 37216 62129 37244
rect 61896 37204 61902 37216
rect 62117 37213 62129 37216
rect 62163 37213 62175 37247
rect 62117 37207 62175 37213
rect 63770 37204 63776 37256
rect 63828 37244 63834 37256
rect 64049 37247 64107 37253
rect 64049 37244 64061 37247
rect 63828 37216 64061 37244
rect 63828 37204 63834 37216
rect 64049 37213 64061 37216
rect 64095 37213 64107 37247
rect 65978 37244 65984 37256
rect 65939 37216 65984 37244
rect 64049 37207 64107 37213
rect 65978 37204 65984 37216
rect 66036 37204 66042 37256
rect 67634 37204 67640 37256
rect 67692 37244 67698 37256
rect 68373 37247 68431 37253
rect 68373 37244 68385 37247
rect 67692 37216 68385 37244
rect 67692 37204 67698 37216
rect 68373 37213 68385 37216
rect 68419 37213 68431 37247
rect 68373 37207 68431 37213
rect 69474 37204 69480 37256
rect 69532 37244 69538 37256
rect 69753 37247 69811 37253
rect 69753 37244 69765 37247
rect 69532 37216 69765 37244
rect 69532 37204 69538 37216
rect 69753 37213 69765 37216
rect 69799 37213 69811 37247
rect 69753 37207 69811 37213
rect 71406 37204 71412 37256
rect 71464 37244 71470 37256
rect 71685 37247 71743 37253
rect 71685 37244 71697 37247
rect 71464 37216 71697 37244
rect 71464 37204 71470 37216
rect 71685 37213 71697 37216
rect 71731 37213 71743 37247
rect 71685 37207 71743 37213
rect 73338 37204 73344 37256
rect 73396 37244 73402 37256
rect 73617 37247 73675 37253
rect 73617 37244 73629 37247
rect 73396 37216 73629 37244
rect 73396 37204 73402 37216
rect 73617 37213 73629 37216
rect 73663 37213 73675 37247
rect 73617 37207 73675 37213
rect 75178 37204 75184 37256
rect 75236 37244 75242 37256
rect 75365 37247 75423 37253
rect 75365 37244 75377 37247
rect 75236 37216 75377 37244
rect 75236 37204 75242 37216
rect 75365 37213 75377 37216
rect 75411 37213 75423 37247
rect 76101 37247 76159 37253
rect 76101 37244 76113 37247
rect 75365 37207 75423 37213
rect 75472 37216 76113 37244
rect 42794 37136 42800 37188
rect 42852 37136 42858 37188
rect 74718 37136 74724 37188
rect 74776 37176 74782 37188
rect 75472 37176 75500 37216
rect 76101 37213 76113 37216
rect 76147 37213 76159 37247
rect 76926 37244 76932 37256
rect 76887 37216 76932 37244
rect 76101 37207 76159 37213
rect 76926 37204 76932 37216
rect 76984 37204 76990 37256
rect 77665 37247 77723 37253
rect 77665 37213 77677 37247
rect 77711 37213 77723 37247
rect 77665 37207 77723 37213
rect 77680 37176 77708 37207
rect 74776 37148 75500 37176
rect 75932 37148 77708 37176
rect 74776 37136 74782 37148
rect 934 37068 940 37120
rect 992 37108 998 37120
rect 1581 37111 1639 37117
rect 1581 37108 1593 37111
rect 992 37080 1593 37108
rect 992 37068 998 37080
rect 1581 37077 1593 37080
rect 1627 37077 1639 37111
rect 1581 37071 1639 37077
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2832 37080 3065 37108
rect 2832 37068 2838 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 3053 37071 3111 37077
rect 4706 37068 4712 37120
rect 4764 37108 4770 37120
rect 4985 37111 5043 37117
rect 4985 37108 4997 37111
rect 4764 37080 4997 37108
rect 4764 37068 4770 37080
rect 4985 37077 4997 37080
rect 5031 37077 5043 37111
rect 4985 37071 5043 37077
rect 6638 37068 6644 37120
rect 6696 37108 6702 37120
rect 6917 37111 6975 37117
rect 6917 37108 6929 37111
rect 6696 37080 6929 37108
rect 6696 37068 6702 37080
rect 6917 37077 6929 37080
rect 6963 37077 6975 37111
rect 6917 37071 6975 37077
rect 8478 37068 8484 37120
rect 8536 37108 8542 37120
rect 9125 37111 9183 37117
rect 9125 37108 9137 37111
rect 8536 37080 9137 37108
rect 8536 37068 8542 37080
rect 9125 37077 9137 37080
rect 9171 37077 9183 37111
rect 9125 37071 9183 37077
rect 10410 37068 10416 37120
rect 10468 37108 10474 37120
rect 10689 37111 10747 37117
rect 10689 37108 10701 37111
rect 10468 37080 10701 37108
rect 10468 37068 10474 37080
rect 10689 37077 10701 37080
rect 10735 37077 10747 37111
rect 10689 37071 10747 37077
rect 12342 37068 12348 37120
rect 12400 37108 12406 37120
rect 12621 37111 12679 37117
rect 12621 37108 12633 37111
rect 12400 37080 12633 37108
rect 12400 37068 12406 37080
rect 12621 37077 12633 37080
rect 12667 37077 12679 37111
rect 12621 37071 12679 37077
rect 14274 37068 14280 37120
rect 14332 37108 14338 37120
rect 14553 37111 14611 37117
rect 14553 37108 14565 37111
rect 14332 37080 14565 37108
rect 14332 37068 14338 37080
rect 14553 37077 14565 37080
rect 14599 37077 14611 37111
rect 14553 37071 14611 37077
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 16853 37111 16911 37117
rect 16853 37108 16865 37111
rect 16632 37080 16865 37108
rect 16632 37068 16638 37080
rect 16853 37077 16865 37080
rect 16899 37077 16911 37111
rect 16853 37071 16911 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18104 37080 18337 37108
rect 18104 37068 18110 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 46566 37068 46572 37120
rect 46624 37108 46630 37120
rect 46753 37111 46811 37117
rect 46753 37108 46765 37111
rect 46624 37080 46765 37108
rect 46624 37068 46630 37080
rect 46753 37077 46765 37080
rect 46799 37077 46811 37111
rect 46753 37071 46811 37077
rect 48593 37111 48651 37117
rect 48593 37077 48605 37111
rect 48639 37108 48651 37111
rect 48866 37108 48872 37120
rect 48639 37080 48872 37108
rect 48639 37077 48651 37080
rect 48593 37071 48651 37077
rect 48866 37068 48872 37080
rect 48924 37068 48930 37120
rect 50525 37111 50583 37117
rect 50525 37077 50537 37111
rect 50571 37108 50583 37111
rect 50798 37108 50804 37120
rect 50571 37080 50804 37108
rect 50571 37077 50583 37080
rect 50525 37071 50583 37077
rect 50798 37068 50804 37080
rect 50856 37068 50862 37120
rect 52454 37068 52460 37120
rect 52512 37108 52518 37120
rect 52733 37111 52791 37117
rect 52733 37108 52745 37111
rect 52512 37080 52745 37108
rect 52512 37068 52518 37080
rect 52733 37077 52745 37080
rect 52779 37077 52791 37111
rect 54386 37108 54392 37120
rect 54347 37080 54392 37108
rect 52733 37071 52791 37077
rect 54386 37068 54392 37080
rect 54444 37068 54450 37120
rect 56042 37068 56048 37120
rect 56100 37108 56106 37120
rect 56229 37111 56287 37117
rect 56229 37108 56241 37111
rect 56100 37080 56241 37108
rect 56100 37068 56106 37080
rect 56229 37077 56241 37080
rect 56275 37077 56287 37111
rect 56229 37071 56287 37077
rect 58161 37111 58219 37117
rect 58161 37077 58173 37111
rect 58207 37108 58219 37111
rect 58434 37108 58440 37120
rect 58207 37080 58440 37108
rect 58207 37077 58219 37080
rect 58161 37071 58219 37077
rect 58434 37068 58440 37080
rect 58492 37068 58498 37120
rect 60461 37111 60519 37117
rect 60461 37077 60473 37111
rect 60507 37108 60519 37111
rect 60642 37108 60648 37120
rect 60507 37080 60648 37108
rect 60507 37077 60519 37080
rect 60461 37071 60519 37077
rect 60642 37068 60648 37080
rect 60700 37068 60706 37120
rect 61930 37108 61936 37120
rect 61891 37080 61936 37108
rect 61930 37068 61936 37080
rect 61988 37068 61994 37120
rect 63862 37108 63868 37120
rect 63823 37080 63868 37108
rect 63862 37068 63868 37080
rect 63920 37068 63926 37120
rect 65797 37111 65855 37117
rect 65797 37077 65809 37111
rect 65843 37108 65855 37111
rect 66162 37108 66168 37120
rect 65843 37080 66168 37108
rect 65843 37077 65855 37080
rect 65797 37071 65855 37077
rect 66162 37068 66168 37080
rect 66220 37068 66226 37120
rect 68186 37108 68192 37120
rect 68147 37080 68192 37108
rect 68186 37068 68192 37080
rect 68244 37068 68250 37120
rect 69566 37108 69572 37120
rect 69527 37080 69572 37108
rect 69566 37068 69572 37080
rect 69624 37068 69630 37120
rect 71498 37108 71504 37120
rect 71459 37080 71504 37108
rect 71498 37068 71504 37080
rect 71556 37068 71562 37120
rect 73433 37111 73491 37117
rect 73433 37077 73445 37111
rect 73479 37108 73491 37111
rect 73706 37108 73712 37120
rect 73479 37080 73712 37108
rect 73479 37077 73491 37080
rect 73433 37071 73491 37077
rect 73706 37068 73712 37080
rect 73764 37068 73770 37120
rect 75086 37068 75092 37120
rect 75144 37108 75150 37120
rect 75932 37117 75960 37148
rect 75181 37111 75239 37117
rect 75181 37108 75193 37111
rect 75144 37080 75193 37108
rect 75144 37068 75150 37080
rect 75181 37077 75193 37080
rect 75227 37077 75239 37111
rect 75181 37071 75239 37077
rect 75917 37111 75975 37117
rect 75917 37077 75929 37111
rect 75963 37077 75975 37111
rect 75917 37071 75975 37077
rect 1104 37018 78844 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 78844 37018
rect 1104 36944 78844 36966
rect 73706 36904 73712 36916
rect 73667 36876 73712 36904
rect 73706 36864 73712 36876
rect 73764 36864 73770 36916
rect 74718 36904 74724 36916
rect 74679 36876 74724 36904
rect 74718 36864 74724 36876
rect 74776 36864 74782 36916
rect 75086 36904 75092 36916
rect 75047 36876 75092 36904
rect 75086 36864 75092 36876
rect 75144 36864 75150 36916
rect 76742 36864 76748 36916
rect 76800 36904 76806 36916
rect 77113 36907 77171 36913
rect 77113 36904 77125 36907
rect 76800 36876 77125 36904
rect 76800 36864 76806 36876
rect 77113 36873 77125 36876
rect 77159 36873 77171 36907
rect 77113 36867 77171 36873
rect 33318 36728 33324 36780
rect 33376 36768 33382 36780
rect 33413 36771 33471 36777
rect 33413 36768 33425 36771
rect 33376 36740 33425 36768
rect 33376 36728 33382 36740
rect 33413 36737 33425 36740
rect 33459 36737 33471 36771
rect 33413 36731 33471 36737
rect 40954 36728 40960 36780
rect 41012 36768 41018 36780
rect 41049 36771 41107 36777
rect 41049 36768 41061 36771
rect 41012 36740 41061 36768
rect 41012 36728 41018 36740
rect 41049 36737 41061 36740
rect 41095 36737 41107 36771
rect 41049 36731 41107 36737
rect 76190 36728 76196 36780
rect 76248 36768 76254 36780
rect 76929 36771 76987 36777
rect 76929 36768 76941 36771
rect 76248 36740 76941 36768
rect 76248 36728 76254 36740
rect 76929 36737 76941 36740
rect 76975 36737 76987 36771
rect 77662 36768 77668 36780
rect 77623 36740 77668 36768
rect 76929 36731 76987 36737
rect 77662 36728 77668 36740
rect 77720 36728 77726 36780
rect 33689 36703 33747 36709
rect 33689 36700 33701 36703
rect 33336 36672 33701 36700
rect 33336 36644 33364 36672
rect 33689 36669 33701 36672
rect 33735 36669 33747 36703
rect 41322 36700 41328 36712
rect 41283 36672 41328 36700
rect 33689 36663 33747 36669
rect 41322 36660 41328 36672
rect 41380 36660 41386 36712
rect 73614 36660 73620 36712
rect 73672 36700 73678 36712
rect 73801 36703 73859 36709
rect 73801 36700 73813 36703
rect 73672 36672 73813 36700
rect 73672 36660 73678 36672
rect 73801 36669 73813 36672
rect 73847 36669 73859 36703
rect 73982 36700 73988 36712
rect 73943 36672 73988 36700
rect 73801 36663 73859 36669
rect 73982 36660 73988 36672
rect 74040 36700 74046 36712
rect 75178 36700 75184 36712
rect 74040 36672 74534 36700
rect 75139 36672 75184 36700
rect 74040 36660 74046 36672
rect 33318 36592 33324 36644
rect 33376 36592 33382 36644
rect 74506 36632 74534 36672
rect 75178 36660 75184 36672
rect 75236 36660 75242 36712
rect 75273 36703 75331 36709
rect 75273 36669 75285 36703
rect 75319 36669 75331 36703
rect 75273 36663 75331 36669
rect 75288 36632 75316 36663
rect 77846 36632 77852 36644
rect 74506 36604 75316 36632
rect 77807 36604 77852 36632
rect 77846 36592 77852 36604
rect 77904 36592 77910 36644
rect 73341 36567 73399 36573
rect 73341 36533 73353 36567
rect 73387 36564 73399 36567
rect 73798 36564 73804 36576
rect 73387 36536 73804 36564
rect 73387 36533 73399 36536
rect 73341 36527 73399 36533
rect 73798 36524 73804 36536
rect 73856 36524 73862 36576
rect 1104 36474 78844 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 78844 36474
rect 1104 36400 78844 36422
rect 73617 36295 73675 36301
rect 73617 36261 73629 36295
rect 73663 36292 73675 36295
rect 73663 36264 74534 36292
rect 73663 36261 73675 36264
rect 73617 36255 73675 36261
rect 74506 36224 74534 36264
rect 77662 36224 77668 36236
rect 74506 36196 77668 36224
rect 77662 36184 77668 36196
rect 77720 36184 77726 36236
rect 73798 36156 73804 36168
rect 73759 36128 73804 36156
rect 73798 36116 73804 36128
rect 73856 36116 73862 36168
rect 77110 36116 77116 36168
rect 77168 36156 77174 36168
rect 77389 36159 77447 36165
rect 77389 36156 77401 36159
rect 77168 36128 77401 36156
rect 77168 36116 77174 36128
rect 77389 36125 77401 36128
rect 77435 36125 77447 36159
rect 77389 36119 77447 36125
rect 77849 36159 77907 36165
rect 77849 36125 77861 36159
rect 77895 36125 77907 36159
rect 77849 36119 77907 36125
rect 73154 36048 73160 36100
rect 73212 36088 73218 36100
rect 77864 36088 77892 36119
rect 73212 36060 77892 36088
rect 73212 36048 73218 36060
rect 76742 35980 76748 36032
rect 76800 36020 76806 36032
rect 77205 36023 77263 36029
rect 77205 36020 77217 36023
rect 76800 35992 77217 36020
rect 76800 35980 76806 35992
rect 77205 35989 77217 35992
rect 77251 35989 77263 36023
rect 78030 36020 78036 36032
rect 77991 35992 78036 36020
rect 77205 35983 77263 35989
rect 78030 35980 78036 35992
rect 78088 35980 78094 36032
rect 1104 35930 78844 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 78844 35930
rect 1104 35856 78844 35878
rect 71498 35816 71504 35828
rect 71459 35788 71504 35816
rect 71498 35776 71504 35788
rect 71556 35776 71562 35828
rect 72329 35819 72387 35825
rect 72329 35785 72341 35819
rect 72375 35816 72387 35819
rect 73154 35816 73160 35828
rect 72375 35788 73160 35816
rect 72375 35785 72387 35788
rect 72329 35779 72387 35785
rect 73154 35776 73160 35788
rect 73212 35776 73218 35828
rect 73246 35748 73252 35760
rect 71700 35720 73252 35748
rect 71406 35572 71412 35624
rect 71464 35612 71470 35624
rect 71700 35621 71728 35720
rect 73246 35708 73252 35720
rect 73304 35748 73310 35760
rect 73982 35748 73988 35760
rect 73304 35720 73988 35748
rect 73304 35708 73310 35720
rect 73982 35708 73988 35720
rect 74040 35708 74046 35760
rect 72513 35683 72571 35689
rect 72513 35649 72525 35683
rect 72559 35649 72571 35683
rect 72513 35643 72571 35649
rect 77941 35683 77999 35689
rect 77941 35649 77953 35683
rect 77987 35680 77999 35683
rect 79042 35680 79048 35692
rect 77987 35652 79048 35680
rect 77987 35649 77999 35652
rect 77941 35643 77999 35649
rect 71593 35615 71651 35621
rect 71593 35612 71605 35615
rect 71464 35584 71605 35612
rect 71464 35572 71470 35584
rect 71593 35581 71605 35584
rect 71639 35581 71651 35615
rect 71593 35575 71651 35581
rect 71685 35615 71743 35621
rect 71685 35581 71697 35615
rect 71731 35581 71743 35615
rect 71685 35575 71743 35581
rect 71133 35547 71191 35553
rect 71133 35513 71145 35547
rect 71179 35544 71191 35547
rect 72528 35544 72556 35643
rect 79042 35640 79048 35652
rect 79100 35640 79106 35692
rect 71179 35516 72556 35544
rect 71179 35513 71191 35516
rect 71133 35507 71191 35513
rect 77754 35476 77760 35488
rect 77715 35448 77760 35476
rect 77754 35436 77760 35448
rect 77812 35436 77818 35488
rect 1104 35386 78844 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 78844 35386
rect 1104 35312 78844 35334
rect 77846 35068 77852 35080
rect 77807 35040 77852 35068
rect 77846 35028 77852 35040
rect 77904 35028 77910 35080
rect 78030 34932 78036 34944
rect 77991 34904 78036 34932
rect 78030 34892 78036 34904
rect 78088 34892 78094 34944
rect 1104 34842 78844 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 78844 34842
rect 1104 34768 78844 34790
rect 69201 34731 69259 34737
rect 69201 34697 69213 34731
rect 69247 34697 69259 34731
rect 69566 34728 69572 34740
rect 69527 34700 69572 34728
rect 69201 34691 69259 34697
rect 69216 34660 69244 34691
rect 69566 34688 69572 34700
rect 69624 34688 69630 34740
rect 70397 34731 70455 34737
rect 70397 34697 70409 34731
rect 70443 34728 70455 34731
rect 70443 34700 74534 34728
rect 70443 34697 70455 34700
rect 70397 34691 70455 34697
rect 74506 34660 74534 34700
rect 76926 34688 76932 34740
rect 76984 34728 76990 34740
rect 77021 34731 77079 34737
rect 77021 34728 77033 34731
rect 76984 34700 77033 34728
rect 76984 34688 76990 34700
rect 77021 34697 77033 34700
rect 77067 34697 77079 34731
rect 77021 34691 77079 34697
rect 77846 34660 77852 34672
rect 69216 34632 70624 34660
rect 74506 34632 77852 34660
rect 69661 34595 69719 34601
rect 69661 34561 69673 34595
rect 69707 34592 69719 34595
rect 69842 34592 69848 34604
rect 69707 34564 69848 34592
rect 69707 34561 69719 34564
rect 69661 34555 69719 34561
rect 69842 34552 69848 34564
rect 69900 34552 69906 34604
rect 70596 34601 70624 34632
rect 77846 34620 77852 34632
rect 77904 34620 77910 34672
rect 70581 34595 70639 34601
rect 70581 34561 70593 34595
rect 70627 34561 70639 34595
rect 77202 34592 77208 34604
rect 77163 34564 77208 34592
rect 70581 34555 70639 34561
rect 77202 34552 77208 34564
rect 77260 34552 77266 34604
rect 77294 34552 77300 34604
rect 77352 34592 77358 34604
rect 77665 34595 77723 34601
rect 77665 34592 77677 34595
rect 77352 34564 77677 34592
rect 77352 34552 77358 34564
rect 77665 34561 77677 34564
rect 77711 34561 77723 34595
rect 77665 34555 77723 34561
rect 69753 34527 69811 34533
rect 69753 34493 69765 34527
rect 69799 34493 69811 34527
rect 69753 34487 69811 34493
rect 68370 34416 68376 34468
rect 68428 34456 68434 34468
rect 69768 34456 69796 34487
rect 73246 34456 73252 34468
rect 68428 34428 73252 34456
rect 68428 34416 68434 34428
rect 73246 34416 73252 34428
rect 73304 34416 73310 34468
rect 77846 34388 77852 34400
rect 77807 34360 77852 34388
rect 77846 34348 77852 34360
rect 77904 34348 77910 34400
rect 1104 34298 78844 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 78844 34298
rect 1104 34224 78844 34246
rect 76190 34184 76196 34196
rect 76151 34156 76196 34184
rect 76190 34144 76196 34156
rect 76248 34144 76254 34196
rect 76837 34187 76895 34193
rect 76837 34153 76849 34187
rect 76883 34184 76895 34187
rect 77202 34184 77208 34196
rect 76883 34156 77208 34184
rect 76883 34153 76895 34156
rect 76837 34147 76895 34153
rect 77202 34144 77208 34156
rect 77260 34144 77266 34196
rect 68370 34048 68376 34060
rect 68331 34020 68376 34048
rect 68370 34008 68376 34020
rect 68428 34008 68434 34060
rect 77110 34008 77116 34060
rect 77168 34048 77174 34060
rect 77389 34051 77447 34057
rect 77389 34048 77401 34051
rect 77168 34020 77401 34048
rect 77168 34008 77174 34020
rect 77389 34017 77401 34020
rect 77435 34017 77447 34051
rect 77389 34011 77447 34017
rect 68097 33983 68155 33989
rect 68097 33949 68109 33983
rect 68143 33980 68155 33983
rect 68186 33980 68192 33992
rect 68143 33952 68192 33980
rect 68143 33949 68155 33952
rect 68097 33943 68155 33949
rect 68186 33940 68192 33952
rect 68244 33940 68250 33992
rect 76377 33983 76435 33989
rect 76377 33949 76389 33983
rect 76423 33980 76435 33983
rect 77202 33980 77208 33992
rect 76423 33952 77208 33980
rect 76423 33949 76435 33952
rect 76377 33943 76435 33949
rect 77202 33940 77208 33952
rect 77260 33940 77266 33992
rect 76926 33872 76932 33924
rect 76984 33912 76990 33924
rect 77297 33915 77355 33921
rect 77297 33912 77309 33915
rect 76984 33884 77309 33912
rect 76984 33872 76990 33884
rect 77297 33881 77309 33884
rect 77343 33881 77355 33915
rect 77297 33875 77355 33881
rect 67726 33844 67732 33856
rect 67687 33816 67732 33844
rect 67726 33804 67732 33816
rect 67784 33804 67790 33856
rect 68189 33847 68247 33853
rect 68189 33813 68201 33847
rect 68235 33844 68247 33847
rect 68370 33844 68376 33856
rect 68235 33816 68376 33844
rect 68235 33813 68247 33816
rect 68189 33807 68247 33813
rect 68370 33804 68376 33816
rect 68428 33804 68434 33856
rect 76742 33804 76748 33856
rect 76800 33844 76806 33856
rect 77205 33847 77263 33853
rect 77205 33844 77217 33847
rect 76800 33816 77217 33844
rect 76800 33804 76806 33816
rect 77205 33813 77217 33816
rect 77251 33813 77263 33847
rect 77205 33807 77263 33813
rect 1104 33754 78844 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 78844 33754
rect 1104 33680 78844 33702
rect 72145 33643 72203 33649
rect 72145 33609 72157 33643
rect 72191 33640 72203 33643
rect 73246 33640 73252 33652
rect 72191 33612 73252 33640
rect 72191 33609 72203 33612
rect 72145 33603 72203 33609
rect 73246 33600 73252 33612
rect 73304 33600 73310 33652
rect 77202 33640 77208 33652
rect 77163 33612 77208 33640
rect 77202 33600 77208 33612
rect 77260 33600 77266 33652
rect 77573 33643 77631 33649
rect 77573 33609 77585 33643
rect 77619 33640 77631 33643
rect 77754 33640 77760 33652
rect 77619 33612 77760 33640
rect 77619 33609 77631 33612
rect 77573 33603 77631 33609
rect 77754 33600 77760 33612
rect 77812 33600 77818 33652
rect 77938 33572 77944 33584
rect 74506 33544 77944 33572
rect 67726 33464 67732 33516
rect 67784 33504 67790 33516
rect 68465 33507 68523 33513
rect 68465 33504 68477 33507
rect 67784 33476 68477 33504
rect 67784 33464 67790 33476
rect 68465 33473 68477 33476
rect 68511 33473 68523 33507
rect 68465 33467 68523 33473
rect 68922 33464 68928 33516
rect 68980 33504 68986 33516
rect 71961 33507 72019 33513
rect 71961 33504 71973 33507
rect 68980 33476 71973 33504
rect 68980 33464 68986 33476
rect 71961 33473 71973 33476
rect 72007 33504 72019 33507
rect 74506 33504 74534 33544
rect 77938 33532 77944 33544
rect 77996 33532 78002 33584
rect 72007 33476 74534 33504
rect 77665 33507 77723 33513
rect 72007 33473 72019 33476
rect 71961 33467 72019 33473
rect 77665 33473 77677 33507
rect 77711 33504 77723 33507
rect 78122 33504 78128 33516
rect 77711 33476 78128 33504
rect 77711 33473 77723 33476
rect 77665 33467 77723 33473
rect 78122 33464 78128 33476
rect 78180 33464 78186 33516
rect 77294 33436 77300 33448
rect 74506 33408 77300 33436
rect 68281 33371 68339 33377
rect 68281 33337 68293 33371
rect 68327 33368 68339 33371
rect 74506 33368 74534 33408
rect 77294 33396 77300 33408
rect 77352 33396 77358 33448
rect 77757 33439 77815 33445
rect 77757 33405 77769 33439
rect 77803 33405 77815 33439
rect 77757 33399 77815 33405
rect 68327 33340 74534 33368
rect 68327 33337 68339 33340
rect 68281 33331 68339 33337
rect 77110 33328 77116 33380
rect 77168 33368 77174 33380
rect 77772 33368 77800 33399
rect 77168 33340 77800 33368
rect 77168 33328 77174 33340
rect 1104 33210 78844 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 78844 33210
rect 1104 33136 78844 33158
rect 78030 33028 78036 33040
rect 77991 33000 78036 33028
rect 78030 32988 78036 33000
rect 78088 32988 78094 33040
rect 76190 32852 76196 32904
rect 76248 32892 76254 32904
rect 77849 32895 77907 32901
rect 77849 32892 77861 32895
rect 76248 32864 77861 32892
rect 76248 32852 76254 32864
rect 77849 32861 77861 32864
rect 77895 32861 77907 32895
rect 77849 32855 77907 32861
rect 1104 32666 78844 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 78844 32666
rect 1104 32592 78844 32614
rect 65978 32416 65984 32428
rect 65939 32388 65984 32416
rect 65978 32376 65984 32388
rect 66036 32376 66042 32428
rect 77662 32416 77668 32428
rect 77623 32388 77668 32416
rect 77662 32376 77668 32388
rect 77720 32376 77726 32428
rect 65797 32215 65855 32221
rect 65797 32181 65809 32215
rect 65843 32212 65855 32215
rect 76190 32212 76196 32224
rect 65843 32184 76196 32212
rect 65843 32181 65855 32184
rect 65797 32175 65855 32181
rect 76190 32172 76196 32184
rect 76248 32172 76254 32224
rect 77846 32212 77852 32224
rect 77807 32184 77852 32212
rect 77846 32172 77852 32184
rect 77904 32172 77910 32224
rect 1104 32122 78844 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 78844 32122
rect 1104 32048 78844 32070
rect 65613 32011 65671 32017
rect 65613 31977 65625 32011
rect 65659 32008 65671 32011
rect 65978 32008 65984 32020
rect 65659 31980 65984 32008
rect 65659 31977 65671 31980
rect 65613 31971 65671 31977
rect 65978 31968 65984 31980
rect 66036 31968 66042 32020
rect 68922 31940 68928 31952
rect 62868 31912 68928 31940
rect 49970 31764 49976 31816
rect 50028 31804 50034 31816
rect 62868 31813 62896 31912
rect 68922 31900 68928 31912
rect 68980 31900 68986 31952
rect 66165 31875 66223 31881
rect 66165 31872 66177 31875
rect 63052 31844 66177 31872
rect 63052 31816 63080 31844
rect 66165 31841 66177 31844
rect 66211 31841 66223 31875
rect 66165 31835 66223 31841
rect 62853 31807 62911 31813
rect 62853 31804 62865 31807
rect 50028 31776 62865 31804
rect 50028 31764 50034 31776
rect 62853 31773 62865 31776
rect 62899 31773 62911 31807
rect 63034 31804 63040 31816
rect 62995 31776 63040 31804
rect 62853 31767 62911 31773
rect 63034 31764 63040 31776
rect 63092 31764 63098 31816
rect 63494 31764 63500 31816
rect 63552 31804 63558 31816
rect 64049 31807 64107 31813
rect 64049 31804 64061 31807
rect 63552 31776 64061 31804
rect 63552 31764 63558 31776
rect 64049 31773 64061 31776
rect 64095 31773 64107 31807
rect 64049 31767 64107 31773
rect 64325 31807 64383 31813
rect 64325 31773 64337 31807
rect 64371 31804 64383 31807
rect 77662 31804 77668 31816
rect 64371 31776 77668 31804
rect 64371 31773 64383 31776
rect 64325 31767 64383 31773
rect 77662 31764 77668 31776
rect 77720 31764 77726 31816
rect 65981 31739 66039 31745
rect 65981 31705 65993 31739
rect 66027 31736 66039 31739
rect 66162 31736 66168 31748
rect 66027 31708 66168 31736
rect 66027 31705 66039 31708
rect 65981 31699 66039 31705
rect 66162 31696 66168 31708
rect 66220 31696 66226 31748
rect 66070 31628 66076 31680
rect 66128 31668 66134 31680
rect 66128 31640 66173 31668
rect 66128 31628 66134 31640
rect 1104 31578 78844 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 78844 31578
rect 1104 31504 78844 31526
rect 61930 31464 61936 31476
rect 61891 31436 61936 31464
rect 61930 31424 61936 31436
rect 61988 31424 61994 31476
rect 63494 31464 63500 31476
rect 63455 31436 63500 31464
rect 63494 31424 63500 31436
rect 63552 31424 63558 31476
rect 63862 31464 63868 31476
rect 63823 31436 63868 31464
rect 63862 31424 63868 31436
rect 63920 31424 63926 31476
rect 63957 31331 64015 31337
rect 63957 31297 63969 31331
rect 64003 31328 64015 31331
rect 64138 31328 64144 31340
rect 64003 31300 64144 31328
rect 64003 31297 64015 31300
rect 63957 31291 64015 31297
rect 64138 31288 64144 31300
rect 64196 31288 64202 31340
rect 77662 31328 77668 31340
rect 77623 31300 77668 31328
rect 77662 31288 77668 31300
rect 77720 31288 77726 31340
rect 61838 31220 61844 31272
rect 61896 31260 61902 31272
rect 62025 31263 62083 31269
rect 62025 31260 62037 31263
rect 61896 31232 62037 31260
rect 61896 31220 61902 31232
rect 62025 31229 62037 31232
rect 62071 31229 62083 31263
rect 62025 31223 62083 31229
rect 62117 31263 62175 31269
rect 62117 31229 62129 31263
rect 62163 31260 62175 31263
rect 63034 31260 63040 31272
rect 62163 31232 63040 31260
rect 62163 31229 62175 31232
rect 62117 31223 62175 31229
rect 61010 31152 61016 31204
rect 61068 31192 61074 31204
rect 62132 31192 62160 31223
rect 63034 31220 63040 31232
rect 63092 31260 63098 31272
rect 64049 31263 64107 31269
rect 64049 31260 64061 31263
rect 63092 31232 64061 31260
rect 63092 31220 63098 31232
rect 64049 31229 64061 31232
rect 64095 31229 64107 31263
rect 64049 31223 64107 31229
rect 61068 31164 62160 31192
rect 61068 31152 61074 31164
rect 61565 31127 61623 31133
rect 61565 31093 61577 31127
rect 61611 31124 61623 31127
rect 62114 31124 62120 31136
rect 61611 31096 62120 31124
rect 61611 31093 61623 31096
rect 61565 31087 61623 31093
rect 62114 31084 62120 31096
rect 62172 31084 62178 31136
rect 77846 31124 77852 31136
rect 77807 31096 77852 31124
rect 77846 31084 77852 31096
rect 77904 31084 77910 31136
rect 1104 31034 78844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 78844 31034
rect 1104 30960 78844 30982
rect 62114 30784 62120 30796
rect 62075 30756 62120 30784
rect 62114 30744 62120 30756
rect 62172 30744 62178 30796
rect 62393 30719 62451 30725
rect 62393 30685 62405 30719
rect 62439 30716 62451 30719
rect 77662 30716 77668 30728
rect 62439 30688 77668 30716
rect 62439 30685 62451 30688
rect 62393 30679 62451 30685
rect 77662 30676 77668 30688
rect 77720 30676 77726 30728
rect 1104 30490 78844 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 78844 30490
rect 1104 30416 78844 30438
rect 58434 30308 58440 30320
rect 58395 30280 58440 30308
rect 58434 30268 58440 30280
rect 58492 30268 58498 30320
rect 77665 30243 77723 30249
rect 77665 30240 77677 30243
rect 64846 30212 77677 30240
rect 58342 30132 58348 30184
rect 58400 30172 58406 30184
rect 58529 30175 58587 30181
rect 58529 30172 58541 30175
rect 58400 30144 58541 30172
rect 58400 30132 58406 30144
rect 58529 30141 58541 30144
rect 58575 30141 58587 30175
rect 58529 30135 58587 30141
rect 58713 30175 58771 30181
rect 58713 30141 58725 30175
rect 58759 30141 58771 30175
rect 58713 30135 58771 30141
rect 60277 30175 60335 30181
rect 60277 30141 60289 30175
rect 60323 30172 60335 30175
rect 60458 30172 60464 30184
rect 60323 30144 60464 30172
rect 60323 30141 60335 30144
rect 60277 30135 60335 30141
rect 58728 30104 58756 30135
rect 60458 30132 60464 30144
rect 60516 30132 60522 30184
rect 60553 30175 60611 30181
rect 60553 30141 60565 30175
rect 60599 30172 60611 30175
rect 64846 30172 64874 30212
rect 77665 30209 77677 30212
rect 77711 30209 77723 30243
rect 77665 30203 77723 30209
rect 60599 30144 64874 30172
rect 60599 30141 60611 30144
rect 60553 30135 60611 30141
rect 61010 30104 61016 30116
rect 58728 30076 61016 30104
rect 61010 30064 61016 30076
rect 61068 30064 61074 30116
rect 77846 30104 77852 30116
rect 77807 30076 77852 30104
rect 77846 30064 77852 30076
rect 77904 30064 77910 30116
rect 58069 30039 58127 30045
rect 58069 30005 58081 30039
rect 58115 30036 58127 30039
rect 58710 30036 58716 30048
rect 58115 30008 58716 30036
rect 58115 30005 58127 30008
rect 58069 29999 58127 30005
rect 58710 29996 58716 30008
rect 58768 29996 58774 30048
rect 1104 29946 78844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 78844 29946
rect 1104 29872 78844 29894
rect 60458 29832 60464 29844
rect 60419 29804 60464 29832
rect 60458 29792 60464 29804
rect 60516 29792 60522 29844
rect 58710 29696 58716 29708
rect 58671 29668 58716 29696
rect 58710 29656 58716 29668
rect 58768 29656 58774 29708
rect 61010 29696 61016 29708
rect 60971 29668 61016 29696
rect 61010 29656 61016 29668
rect 61068 29656 61074 29708
rect 58989 29631 59047 29637
rect 58989 29597 59001 29631
rect 59035 29628 59047 29631
rect 77849 29631 77907 29637
rect 77849 29628 77861 29631
rect 59035 29600 77861 29628
rect 59035 29597 59047 29600
rect 58989 29591 59047 29597
rect 77849 29597 77861 29600
rect 77895 29597 77907 29631
rect 77849 29591 77907 29597
rect 60642 29520 60648 29572
rect 60700 29560 60706 29572
rect 60829 29563 60887 29569
rect 60829 29560 60841 29563
rect 60700 29532 60841 29560
rect 60700 29520 60706 29532
rect 60829 29529 60841 29532
rect 60875 29529 60887 29563
rect 60829 29523 60887 29529
rect 60734 29452 60740 29504
rect 60792 29492 60798 29504
rect 60921 29495 60979 29501
rect 60921 29492 60933 29495
rect 60792 29464 60933 29492
rect 60792 29452 60798 29464
rect 60921 29461 60933 29464
rect 60967 29461 60979 29495
rect 78030 29492 78036 29504
rect 77991 29464 78036 29492
rect 60921 29455 60979 29461
rect 78030 29452 78036 29464
rect 78088 29452 78094 29504
rect 1104 29402 78844 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 78844 29402
rect 1104 29328 78844 29350
rect 1104 28858 78844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 78844 28858
rect 1104 28784 78844 28806
rect 77846 28540 77852 28552
rect 77807 28512 77852 28540
rect 77846 28500 77852 28512
rect 77904 28500 77910 28552
rect 78030 28404 78036 28416
rect 77991 28376 78036 28404
rect 78030 28364 78036 28376
rect 78088 28364 78094 28416
rect 1104 28314 78844 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 78844 28314
rect 1104 28240 78844 28262
rect 56318 28064 56324 28076
rect 56279 28036 56324 28064
rect 56318 28024 56324 28036
rect 56376 28024 56382 28076
rect 56413 27863 56471 27869
rect 56413 27829 56425 27863
rect 56459 27860 56471 27863
rect 77846 27860 77852 27872
rect 56459 27832 77852 27860
rect 56459 27829 56471 27832
rect 56413 27823 56471 27829
rect 77846 27820 77852 27832
rect 77904 27820 77910 27872
rect 1104 27770 78844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 78844 27770
rect 1104 27696 78844 27718
rect 55677 27659 55735 27665
rect 55677 27625 55689 27659
rect 55723 27656 55735 27659
rect 56318 27656 56324 27668
rect 55723 27628 56324 27656
rect 55723 27625 55735 27628
rect 55677 27619 55735 27625
rect 56318 27616 56324 27628
rect 56376 27616 56382 27668
rect 52638 27480 52644 27532
rect 52696 27520 52702 27532
rect 54573 27523 54631 27529
rect 54573 27520 54585 27523
rect 52696 27492 54585 27520
rect 52696 27480 52702 27492
rect 54573 27489 54585 27492
rect 54619 27520 54631 27523
rect 56229 27523 56287 27529
rect 56229 27520 56241 27523
rect 54619 27492 56241 27520
rect 54619 27489 54631 27492
rect 54573 27483 54631 27489
rect 56229 27489 56241 27492
rect 56275 27489 56287 27523
rect 56229 27483 56287 27489
rect 54386 27452 54392 27464
rect 54347 27424 54392 27452
rect 54386 27412 54392 27424
rect 54444 27412 54450 27464
rect 56042 27452 56048 27464
rect 56003 27424 56048 27452
rect 56042 27412 56048 27424
rect 56100 27412 56106 27464
rect 76190 27412 76196 27464
rect 76248 27452 76254 27464
rect 77849 27455 77907 27461
rect 77849 27452 77861 27455
rect 76248 27424 77861 27452
rect 76248 27412 76254 27424
rect 77849 27421 77861 27424
rect 77895 27421 77907 27455
rect 77849 27415 77907 27421
rect 54018 27316 54024 27328
rect 53979 27288 54024 27316
rect 54018 27276 54024 27288
rect 54076 27276 54082 27328
rect 54481 27319 54539 27325
rect 54481 27285 54493 27319
rect 54527 27316 54539 27319
rect 54570 27316 54576 27328
rect 54527 27288 54576 27316
rect 54527 27285 54539 27288
rect 54481 27279 54539 27285
rect 54570 27276 54576 27288
rect 54628 27276 54634 27328
rect 56137 27319 56195 27325
rect 56137 27285 56149 27319
rect 56183 27316 56195 27319
rect 56410 27316 56416 27328
rect 56183 27288 56416 27316
rect 56183 27285 56195 27288
rect 56137 27279 56195 27285
rect 56410 27276 56416 27288
rect 56468 27276 56474 27328
rect 78030 27316 78036 27328
rect 77991 27288 78036 27316
rect 78030 27276 78036 27288
rect 78088 27276 78094 27328
rect 1104 27226 78844 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 78844 27226
rect 1104 27152 78844 27174
rect 54018 27004 54024 27056
rect 54076 27044 54082 27056
rect 54665 27047 54723 27053
rect 54665 27044 54677 27047
rect 54076 27016 54677 27044
rect 54076 27004 54082 27016
rect 54665 27013 54677 27016
rect 54711 27013 54723 27047
rect 54665 27007 54723 27013
rect 77662 26976 77668 26988
rect 77623 26948 77668 26976
rect 77662 26936 77668 26948
rect 77720 26936 77726 26988
rect 54757 26775 54815 26781
rect 54757 26741 54769 26775
rect 54803 26772 54815 26775
rect 76190 26772 76196 26784
rect 54803 26744 76196 26772
rect 54803 26741 54815 26744
rect 54757 26735 54815 26741
rect 76190 26732 76196 26744
rect 76248 26732 76254 26784
rect 77846 26772 77852 26784
rect 77807 26744 77852 26772
rect 77846 26732 77852 26744
rect 77904 26732 77910 26784
rect 1104 26682 78844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 78844 26682
rect 1104 26608 78844 26630
rect 52089 26503 52147 26509
rect 52089 26469 52101 26503
rect 52135 26500 52147 26503
rect 52135 26472 53420 26500
rect 52135 26469 52147 26472
rect 52089 26463 52147 26469
rect 50706 26392 50712 26444
rect 50764 26432 50770 26444
rect 52638 26432 52644 26444
rect 50764 26404 52644 26432
rect 50764 26392 50770 26404
rect 52638 26392 52644 26404
rect 52696 26392 52702 26444
rect 52454 26364 52460 26376
rect 52415 26336 52460 26364
rect 52454 26324 52460 26336
rect 52512 26324 52518 26376
rect 53392 26373 53420 26472
rect 53377 26367 53435 26373
rect 53377 26333 53389 26367
rect 53423 26333 53435 26367
rect 53377 26327 53435 26333
rect 52549 26299 52607 26305
rect 52549 26265 52561 26299
rect 52595 26296 52607 26299
rect 52914 26296 52920 26308
rect 52595 26268 52920 26296
rect 52595 26265 52607 26268
rect 52549 26259 52607 26265
rect 52914 26256 52920 26268
rect 52972 26256 52978 26308
rect 53561 26299 53619 26305
rect 53561 26265 53573 26299
rect 53607 26296 53619 26299
rect 77662 26296 77668 26308
rect 53607 26268 77668 26296
rect 53607 26265 53619 26268
rect 53561 26259 53619 26265
rect 77662 26256 77668 26268
rect 77720 26256 77726 26308
rect 1104 26138 78844 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 78844 26138
rect 1104 26064 78844 26086
rect 77662 25888 77668 25900
rect 77623 25860 77668 25888
rect 77662 25848 77668 25860
rect 77720 25848 77726 25900
rect 77846 25684 77852 25696
rect 77807 25656 77852 25684
rect 77846 25644 77852 25656
rect 77904 25644 77910 25696
rect 1104 25594 78844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 78844 25594
rect 1104 25520 78844 25542
rect 50706 25344 50712 25356
rect 50667 25316 50712 25344
rect 50706 25304 50712 25316
rect 50764 25304 50770 25356
rect 50525 25279 50583 25285
rect 50525 25245 50537 25279
rect 50571 25276 50583 25279
rect 50798 25276 50804 25288
rect 50571 25248 50804 25276
rect 50571 25245 50583 25248
rect 50525 25239 50583 25245
rect 50798 25236 50804 25248
rect 50856 25236 50862 25288
rect 51445 25211 51503 25217
rect 51445 25208 51457 25211
rect 50172 25180 51457 25208
rect 50172 25149 50200 25180
rect 51445 25177 51457 25180
rect 51491 25177 51503 25211
rect 51445 25171 51503 25177
rect 50157 25143 50215 25149
rect 50157 25109 50169 25143
rect 50203 25109 50215 25143
rect 50157 25103 50215 25109
rect 50617 25143 50675 25149
rect 50617 25109 50629 25143
rect 50663 25140 50675 25143
rect 50706 25140 50712 25152
rect 50663 25112 50712 25140
rect 50663 25109 50675 25112
rect 50617 25103 50675 25109
rect 50706 25100 50712 25112
rect 50764 25100 50770 25152
rect 51537 25143 51595 25149
rect 51537 25109 51549 25143
rect 51583 25140 51595 25143
rect 77662 25140 77668 25152
rect 51583 25112 77668 25140
rect 51583 25109 51595 25112
rect 51537 25103 51595 25109
rect 77662 25100 77668 25112
rect 77720 25100 77726 25152
rect 1104 25050 78844 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 78844 25050
rect 1104 24976 78844 24998
rect 48866 24936 48872 24948
rect 48827 24908 48872 24936
rect 48866 24896 48872 24908
rect 48924 24896 48930 24948
rect 48961 24803 49019 24809
rect 48961 24769 48973 24803
rect 49007 24800 49019 24803
rect 49142 24800 49148 24812
rect 49007 24772 49148 24800
rect 49007 24769 49019 24772
rect 48961 24763 49019 24769
rect 49142 24760 49148 24772
rect 49200 24760 49206 24812
rect 77662 24800 77668 24812
rect 77623 24772 77668 24800
rect 77662 24760 77668 24772
rect 77720 24760 77726 24812
rect 49053 24735 49111 24741
rect 49053 24701 49065 24735
rect 49099 24732 49111 24735
rect 49694 24732 49700 24744
rect 49099 24704 49700 24732
rect 49099 24701 49111 24704
rect 49053 24695 49111 24701
rect 49694 24692 49700 24704
rect 49752 24732 49758 24744
rect 50614 24732 50620 24744
rect 49752 24704 50620 24732
rect 49752 24692 49758 24704
rect 50614 24692 50620 24704
rect 50672 24692 50678 24744
rect 48501 24599 48559 24605
rect 48501 24565 48513 24599
rect 48547 24596 48559 24599
rect 49234 24596 49240 24608
rect 48547 24568 49240 24596
rect 48547 24565 48559 24568
rect 48501 24559 48559 24565
rect 49234 24556 49240 24568
rect 49292 24556 49298 24608
rect 77846 24596 77852 24608
rect 77807 24568 77852 24596
rect 77846 24556 77852 24568
rect 77904 24556 77910 24608
rect 1104 24506 78844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 78844 24506
rect 1104 24432 78844 24454
rect 49234 24188 49240 24200
rect 49195 24160 49240 24188
rect 49234 24148 49240 24160
rect 49292 24148 49298 24200
rect 49329 24055 49387 24061
rect 49329 24021 49341 24055
rect 49375 24052 49387 24055
rect 77662 24052 77668 24064
rect 49375 24024 77668 24052
rect 49375 24021 49387 24024
rect 49329 24015 49387 24021
rect 77662 24012 77668 24024
rect 77720 24012 77726 24064
rect 1104 23962 78844 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 78844 23962
rect 1104 23888 78844 23910
rect 49694 23848 49700 23860
rect 49655 23820 49700 23848
rect 49694 23808 49700 23820
rect 49752 23808 49758 23860
rect 49602 23712 49608 23724
rect 49563 23684 49608 23712
rect 49602 23672 49608 23684
rect 49660 23672 49666 23724
rect 77297 23715 77355 23721
rect 77297 23712 77309 23715
rect 55186 23684 77309 23712
rect 47026 23604 47032 23656
rect 47084 23644 47090 23656
rect 55186 23644 55214 23684
rect 77297 23681 77309 23684
rect 77343 23712 77355 23715
rect 77665 23715 77723 23721
rect 77665 23712 77677 23715
rect 77343 23684 77677 23712
rect 77343 23681 77355 23684
rect 77297 23675 77355 23681
rect 77665 23681 77677 23684
rect 77711 23681 77723 23715
rect 77665 23675 77723 23681
rect 47084 23616 55214 23644
rect 47084 23604 47090 23616
rect 77846 23576 77852 23588
rect 77807 23548 77852 23576
rect 77846 23536 77852 23548
rect 77904 23536 77910 23588
rect 1104 23418 78844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 78844 23418
rect 1104 23344 78844 23366
rect 47026 23236 47032 23248
rect 46987 23208 47032 23236
rect 47026 23196 47032 23208
rect 47084 23196 47090 23248
rect 77849 23103 77907 23109
rect 77849 23100 77861 23103
rect 77496 23072 77861 23100
rect 46198 22992 46204 23044
rect 46256 23032 46262 23044
rect 46845 23035 46903 23041
rect 46845 23032 46857 23035
rect 46256 23004 46857 23032
rect 46256 22992 46262 23004
rect 46845 23001 46857 23004
rect 46891 23001 46903 23035
rect 46845 22995 46903 23001
rect 77496 22976 77524 23072
rect 77849 23069 77861 23072
rect 77895 23069 77907 23103
rect 77849 23063 77907 23069
rect 77478 22964 77484 22976
rect 77439 22936 77484 22964
rect 77478 22924 77484 22936
rect 77536 22924 77542 22976
rect 78030 22964 78036 22976
rect 77991 22936 78036 22964
rect 78030 22924 78036 22936
rect 78088 22924 78094 22976
rect 1104 22874 78844 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 78844 22874
rect 1104 22800 78844 22822
rect 44818 22760 44824 22772
rect 44779 22732 44824 22760
rect 44818 22720 44824 22732
rect 44876 22720 44882 22772
rect 46198 22760 46204 22772
rect 46159 22732 46204 22760
rect 46198 22720 46204 22732
rect 46256 22720 46262 22772
rect 46566 22760 46572 22772
rect 46527 22732 46572 22760
rect 46566 22720 46572 22732
rect 46624 22720 46630 22772
rect 77478 22760 77484 22772
rect 55186 22732 77484 22760
rect 45186 22652 45192 22704
rect 45244 22692 45250 22704
rect 55186 22692 55214 22732
rect 77478 22720 77484 22732
rect 77536 22720 77542 22772
rect 45244 22664 55214 22692
rect 45244 22652 45250 22664
rect 44913 22627 44971 22633
rect 44913 22593 44925 22627
rect 44959 22624 44971 22627
rect 45278 22624 45284 22636
rect 44959 22596 45284 22624
rect 44959 22593 44971 22596
rect 44913 22587 44971 22593
rect 45278 22584 45284 22596
rect 45336 22584 45342 22636
rect 49970 22624 49976 22636
rect 49931 22596 49976 22624
rect 49970 22584 49976 22596
rect 50028 22584 50034 22636
rect 45005 22559 45063 22565
rect 45005 22525 45017 22559
rect 45051 22525 45063 22559
rect 46658 22556 46664 22568
rect 46619 22528 46664 22556
rect 45005 22519 45063 22525
rect 43162 22448 43168 22500
rect 43220 22488 43226 22500
rect 45020 22488 45048 22519
rect 46658 22516 46664 22528
rect 46716 22516 46722 22568
rect 46753 22559 46811 22565
rect 46753 22525 46765 22559
rect 46799 22525 46811 22559
rect 46753 22519 46811 22525
rect 46768 22488 46796 22519
rect 43220 22460 46796 22488
rect 43220 22448 43226 22460
rect 44453 22423 44511 22429
rect 44453 22389 44465 22423
rect 44499 22420 44511 22423
rect 45002 22420 45008 22432
rect 44499 22392 45008 22420
rect 44499 22389 44511 22392
rect 44453 22383 44511 22389
rect 45002 22380 45008 22392
rect 45060 22380 45066 22432
rect 49602 22380 49608 22432
rect 49660 22420 49666 22432
rect 50065 22423 50123 22429
rect 50065 22420 50077 22423
rect 49660 22392 50077 22420
rect 49660 22380 49666 22392
rect 50065 22389 50077 22392
rect 50111 22389 50123 22423
rect 50065 22383 50123 22389
rect 1104 22330 78844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 78844 22330
rect 1104 22256 78844 22278
rect 45186 22216 45192 22228
rect 45147 22188 45192 22216
rect 45186 22176 45192 22188
rect 45244 22176 45250 22228
rect 41690 22108 41696 22160
rect 41748 22148 41754 22160
rect 43162 22148 43168 22160
rect 41748 22120 43168 22148
rect 41748 22108 41754 22120
rect 43162 22108 43168 22120
rect 43220 22108 43226 22160
rect 40405 22083 40463 22089
rect 40405 22049 40417 22083
rect 40451 22080 40463 22083
rect 41708 22080 41736 22108
rect 43073 22083 43131 22089
rect 40451 22052 41736 22080
rect 41800 22052 43024 22080
rect 40451 22049 40463 22052
rect 40405 22043 40463 22049
rect 36538 21972 36544 22024
rect 36596 22012 36602 22024
rect 40221 22015 40279 22021
rect 40221 22012 40233 22015
rect 36596 21984 40233 22012
rect 36596 21972 36602 21984
rect 40221 21981 40233 21984
rect 40267 22012 40279 22015
rect 41800 22012 41828 22052
rect 40267 21984 41828 22012
rect 40267 21981 40279 21984
rect 40221 21975 40279 21981
rect 42794 21972 42800 22024
rect 42852 22012 42858 22024
rect 42889 22015 42947 22021
rect 42889 22012 42901 22015
rect 42852 21984 42901 22012
rect 42852 21972 42858 21984
rect 42889 21981 42901 21984
rect 42935 21981 42947 22015
rect 42996 22012 43024 22052
rect 43073 22049 43085 22083
rect 43119 22080 43131 22083
rect 43180 22080 43208 22108
rect 49602 22080 49608 22092
rect 43119 22052 43208 22080
rect 43272 22052 49608 22080
rect 43119 22049 43131 22052
rect 43073 22043 43131 22049
rect 43272 22012 43300 22052
rect 49602 22040 49608 22052
rect 49660 22040 49666 22092
rect 42996 21984 43300 22012
rect 43717 22015 43775 22021
rect 42889 21975 42947 21981
rect 43717 21981 43729 22015
rect 43763 21981 43775 22015
rect 45002 22012 45008 22024
rect 44963 21984 45008 22012
rect 43717 21975 43775 21981
rect 43732 21944 43760 21975
rect 45002 21972 45008 21984
rect 45060 21972 45066 22024
rect 77846 22012 77852 22024
rect 77807 21984 77852 22012
rect 77846 21972 77852 21984
rect 77904 21972 77910 22024
rect 42536 21916 43760 21944
rect 42536 21885 42564 21916
rect 42521 21879 42579 21885
rect 42521 21845 42533 21879
rect 42567 21845 42579 21879
rect 42521 21839 42579 21845
rect 42981 21879 43039 21885
rect 42981 21845 42993 21879
rect 43027 21876 43039 21879
rect 43162 21876 43168 21888
rect 43027 21848 43168 21876
rect 43027 21845 43039 21848
rect 42981 21839 43039 21845
rect 43162 21836 43168 21848
rect 43220 21836 43226 21888
rect 43898 21876 43904 21888
rect 43859 21848 43904 21876
rect 43898 21836 43904 21848
rect 43956 21836 43962 21888
rect 78030 21876 78036 21888
rect 77991 21848 78036 21876
rect 78030 21836 78036 21848
rect 78088 21836 78094 21888
rect 1104 21786 78844 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 78844 21786
rect 1104 21712 78844 21734
rect 43898 21632 43904 21684
rect 43956 21672 43962 21684
rect 77846 21672 77852 21684
rect 43956 21644 77852 21672
rect 43956 21632 43962 21644
rect 77846 21632 77852 21644
rect 77904 21632 77910 21684
rect 1104 21242 78844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 78844 21242
rect 1104 21168 78844 21190
rect 40497 20995 40555 21001
rect 40497 20961 40509 20995
rect 40543 20992 40555 20995
rect 41690 20992 41696 21004
rect 40543 20964 41696 20992
rect 40543 20961 40555 20964
rect 40497 20955 40555 20961
rect 41690 20952 41696 20964
rect 41748 20952 41754 21004
rect 40218 20924 40224 20936
rect 40179 20896 40224 20924
rect 40218 20884 40224 20896
rect 40276 20884 40282 20936
rect 41322 20884 41328 20936
rect 41380 20924 41386 20936
rect 41417 20927 41475 20933
rect 41417 20924 41429 20927
rect 41380 20896 41429 20924
rect 41380 20884 41386 20896
rect 41417 20893 41429 20896
rect 41463 20893 41475 20927
rect 77849 20927 77907 20933
rect 77849 20924 77861 20927
rect 41417 20887 41475 20893
rect 77496 20896 77861 20924
rect 41598 20816 41604 20868
rect 41656 20856 41662 20868
rect 77496 20865 77524 20896
rect 77849 20893 77861 20896
rect 77895 20893 77907 20927
rect 77849 20887 77907 20893
rect 77481 20859 77539 20865
rect 77481 20856 77493 20859
rect 41656 20828 77493 20856
rect 41656 20816 41662 20828
rect 77481 20825 77493 20828
rect 77527 20825 77539 20859
rect 77481 20819 77539 20825
rect 39666 20748 39672 20800
rect 39724 20788 39730 20800
rect 39853 20791 39911 20797
rect 39853 20788 39865 20791
rect 39724 20760 39865 20788
rect 39724 20748 39730 20760
rect 39853 20757 39865 20760
rect 39899 20757 39911 20791
rect 39853 20751 39911 20757
rect 40126 20748 40132 20800
rect 40184 20788 40190 20800
rect 40313 20791 40371 20797
rect 40313 20788 40325 20791
rect 40184 20760 40325 20788
rect 40184 20748 40190 20760
rect 40313 20757 40325 20760
rect 40359 20757 40371 20791
rect 40313 20751 40371 20757
rect 41049 20791 41107 20797
rect 41049 20757 41061 20791
rect 41095 20788 41107 20791
rect 41230 20788 41236 20800
rect 41095 20760 41236 20788
rect 41095 20757 41107 20760
rect 41049 20751 41107 20757
rect 41230 20748 41236 20760
rect 41288 20748 41294 20800
rect 41506 20748 41512 20800
rect 41564 20788 41570 20800
rect 78030 20788 78036 20800
rect 41564 20760 41609 20788
rect 77991 20760 78036 20788
rect 41564 20748 41570 20760
rect 78030 20748 78036 20760
rect 78088 20748 78094 20800
rect 1104 20698 78844 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 78844 20698
rect 1104 20624 78844 20646
rect 41417 20587 41475 20593
rect 41417 20553 41429 20587
rect 41463 20584 41475 20587
rect 41598 20584 41604 20596
rect 41463 20556 41604 20584
rect 41463 20553 41475 20556
rect 41417 20547 41475 20553
rect 41598 20544 41604 20556
rect 41656 20544 41662 20596
rect 39666 20448 39672 20460
rect 39627 20420 39672 20448
rect 39666 20408 39672 20420
rect 39724 20408 39730 20460
rect 41230 20448 41236 20460
rect 41191 20420 41236 20448
rect 41230 20408 41236 20420
rect 41288 20408 41294 20460
rect 49970 20408 49976 20460
rect 50028 20448 50034 20460
rect 50341 20451 50399 20457
rect 50341 20448 50353 20451
rect 50028 20420 50353 20448
rect 50028 20408 50034 20420
rect 50341 20417 50353 20420
rect 50387 20417 50399 20451
rect 50341 20411 50399 20417
rect 77665 20451 77723 20457
rect 77665 20417 77677 20451
rect 77711 20417 77723 20451
rect 77665 20411 77723 20417
rect 50982 20380 50988 20392
rect 50943 20352 50988 20380
rect 50982 20340 50988 20352
rect 51040 20380 51046 20392
rect 77110 20380 77116 20392
rect 51040 20352 77116 20380
rect 51040 20340 51046 20352
rect 77110 20340 77116 20352
rect 77168 20340 77174 20392
rect 39853 20315 39911 20321
rect 39853 20281 39865 20315
rect 39899 20312 39911 20315
rect 77680 20312 77708 20411
rect 39899 20284 77708 20312
rect 39899 20281 39911 20284
rect 39853 20275 39911 20281
rect 77846 20244 77852 20256
rect 77807 20216 77852 20244
rect 77846 20204 77852 20216
rect 77904 20204 77910 20256
rect 1104 20154 78844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 78844 20154
rect 1104 20080 78844 20102
rect 1104 19610 78844 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 78844 19610
rect 1104 19536 78844 19558
rect 77294 19320 77300 19372
rect 77352 19360 77358 19372
rect 77665 19363 77723 19369
rect 77665 19360 77677 19363
rect 77352 19332 77677 19360
rect 77352 19320 77358 19332
rect 77665 19329 77677 19332
rect 77711 19329 77723 19363
rect 77665 19323 77723 19329
rect 77294 19156 77300 19168
rect 77255 19128 77300 19156
rect 77294 19116 77300 19128
rect 77352 19116 77358 19168
rect 77846 19156 77852 19168
rect 77807 19128 77852 19156
rect 77846 19116 77852 19128
rect 77904 19116 77910 19168
rect 1104 19066 78844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 78844 19066
rect 1104 18992 78844 19014
rect 37185 18751 37243 18757
rect 37185 18717 37197 18751
rect 37231 18748 37243 18751
rect 37274 18748 37280 18760
rect 37231 18720 37280 18748
rect 37231 18717 37243 18720
rect 37185 18711 37243 18717
rect 37274 18708 37280 18720
rect 37332 18708 37338 18760
rect 37369 18615 37427 18621
rect 37369 18581 37381 18615
rect 37415 18612 37427 18615
rect 77294 18612 77300 18624
rect 37415 18584 77300 18612
rect 37415 18581 37427 18584
rect 37369 18575 37427 18581
rect 77294 18572 77300 18584
rect 77352 18572 77358 18624
rect 1104 18522 78844 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 78844 18522
rect 1104 18448 78844 18470
rect 37274 18408 37280 18420
rect 37235 18380 37280 18408
rect 37274 18368 37280 18380
rect 37332 18368 37338 18420
rect 37642 18408 37648 18420
rect 37603 18380 37648 18408
rect 37642 18368 37648 18380
rect 37700 18368 37706 18420
rect 36262 18232 36268 18284
rect 36320 18272 36326 18284
rect 77297 18275 77355 18281
rect 77297 18272 77309 18275
rect 36320 18244 77309 18272
rect 36320 18232 36326 18244
rect 77297 18241 77309 18244
rect 77343 18272 77355 18275
rect 77665 18275 77723 18281
rect 77665 18272 77677 18275
rect 77343 18244 77677 18272
rect 77343 18241 77355 18244
rect 77297 18235 77355 18241
rect 77665 18241 77677 18244
rect 77711 18241 77723 18275
rect 77665 18235 77723 18241
rect 37550 18164 37556 18216
rect 37608 18204 37614 18216
rect 37737 18207 37795 18213
rect 37737 18204 37749 18207
rect 37608 18176 37749 18204
rect 37608 18164 37614 18176
rect 37737 18173 37749 18176
rect 37783 18173 37795 18207
rect 37737 18167 37795 18173
rect 37829 18207 37887 18213
rect 37829 18173 37841 18207
rect 37875 18173 37887 18207
rect 37829 18167 37887 18173
rect 36722 18096 36728 18148
rect 36780 18136 36786 18148
rect 37844 18136 37872 18167
rect 36780 18108 37872 18136
rect 36780 18096 36786 18108
rect 77846 18068 77852 18080
rect 77807 18040 77852 18068
rect 77846 18028 77852 18040
rect 77904 18028 77910 18080
rect 1104 17978 78844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 78844 17978
rect 1104 17904 78844 17926
rect 36262 17864 36268 17876
rect 36223 17836 36268 17864
rect 36262 17824 36268 17836
rect 36320 17824 36326 17876
rect 34885 17799 34943 17805
rect 34885 17765 34897 17799
rect 34931 17796 34943 17799
rect 34931 17768 36124 17796
rect 34931 17765 34943 17768
rect 34885 17759 34943 17765
rect 33686 17688 33692 17740
rect 33744 17728 33750 17740
rect 35437 17731 35495 17737
rect 35437 17728 35449 17731
rect 33744 17700 35449 17728
rect 33744 17688 33750 17700
rect 35437 17697 35449 17700
rect 35483 17728 35495 17731
rect 35483 17700 35894 17728
rect 35483 17697 35495 17700
rect 35437 17691 35495 17697
rect 35253 17595 35311 17601
rect 35253 17561 35265 17595
rect 35299 17592 35311 17595
rect 35434 17592 35440 17604
rect 35299 17564 35440 17592
rect 35299 17561 35311 17564
rect 35253 17555 35311 17561
rect 35434 17552 35440 17564
rect 35492 17552 35498 17604
rect 35866 17592 35894 17700
rect 36096 17669 36124 17768
rect 36081 17663 36139 17669
rect 36081 17629 36093 17663
rect 36127 17629 36139 17663
rect 77846 17660 77852 17672
rect 77807 17632 77852 17660
rect 36081 17623 36139 17629
rect 77846 17620 77852 17632
rect 77904 17620 77910 17672
rect 36722 17592 36728 17604
rect 35866 17564 36728 17592
rect 36722 17552 36728 17564
rect 36780 17552 36786 17604
rect 35345 17527 35403 17533
rect 35345 17493 35357 17527
rect 35391 17524 35403 17527
rect 35526 17524 35532 17536
rect 35391 17496 35532 17524
rect 35391 17493 35403 17496
rect 35345 17487 35403 17493
rect 35526 17484 35532 17496
rect 35584 17484 35590 17536
rect 78030 17524 78036 17536
rect 77991 17496 78036 17524
rect 78030 17484 78036 17496
rect 78088 17484 78094 17536
rect 1104 17434 78844 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 78844 17434
rect 1104 17360 78844 17382
rect 33318 17280 33324 17332
rect 33376 17320 33382 17332
rect 33413 17323 33471 17329
rect 33413 17320 33425 17323
rect 33376 17292 33425 17320
rect 33376 17280 33382 17292
rect 33413 17289 33425 17292
rect 33459 17289 33471 17323
rect 33413 17283 33471 17289
rect 31662 17212 31668 17264
rect 31720 17252 31726 17264
rect 33686 17252 33692 17264
rect 31720 17224 33692 17252
rect 31720 17212 31726 17224
rect 33686 17212 33692 17224
rect 33744 17212 33750 17264
rect 36538 17252 36544 17264
rect 36499 17224 36544 17252
rect 36538 17212 36544 17224
rect 36596 17212 36602 17264
rect 36722 17252 36728 17264
rect 36683 17224 36728 17252
rect 36722 17212 36728 17224
rect 36780 17212 36786 17264
rect 33502 17116 33508 17128
rect 33463 17088 33508 17116
rect 33502 17076 33508 17088
rect 33560 17076 33566 17128
rect 33704 17125 33732 17212
rect 34241 17187 34299 17193
rect 34241 17153 34253 17187
rect 34287 17153 34299 17187
rect 34241 17147 34299 17153
rect 33689 17119 33747 17125
rect 33689 17085 33701 17119
rect 33735 17085 33747 17119
rect 33689 17079 33747 17085
rect 33045 17051 33103 17057
rect 33045 17017 33057 17051
rect 33091 17048 33103 17051
rect 34256 17048 34284 17147
rect 33091 17020 34284 17048
rect 34425 17051 34483 17057
rect 33091 17017 33103 17020
rect 33045 17011 33103 17017
rect 34425 17017 34437 17051
rect 34471 17048 34483 17051
rect 34471 17020 45554 17048
rect 34471 17017 34483 17020
rect 34425 17011 34483 17017
rect 45526 16980 45554 17020
rect 77846 16980 77852 16992
rect 45526 16952 77852 16980
rect 77846 16940 77852 16952
rect 77904 16940 77910 16992
rect 1104 16890 78844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 78844 16890
rect 1104 16816 78844 16838
rect 31570 16640 31576 16652
rect 31531 16612 31576 16640
rect 31570 16600 31576 16612
rect 31628 16600 31634 16652
rect 31662 16600 31668 16652
rect 31720 16640 31726 16652
rect 31720 16612 31765 16640
rect 31720 16600 31726 16612
rect 31481 16575 31539 16581
rect 31481 16541 31493 16575
rect 31527 16572 31539 16575
rect 32398 16572 32404 16584
rect 31527 16544 32404 16572
rect 31527 16541 31539 16544
rect 31481 16535 31539 16541
rect 32398 16532 32404 16544
rect 32456 16532 32462 16584
rect 77846 16572 77852 16584
rect 77807 16544 77852 16572
rect 77846 16532 77852 16544
rect 77904 16532 77910 16584
rect 31110 16436 31116 16448
rect 31071 16408 31116 16436
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 78030 16436 78036 16448
rect 77991 16408 78036 16436
rect 78030 16396 78036 16408
rect 78088 16396 78094 16448
rect 1104 16346 78844 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 78844 16346
rect 1104 16272 78844 16294
rect 29914 16232 29920 16244
rect 29875 16204 29920 16232
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 31110 16124 31116 16176
rect 31168 16164 31174 16176
rect 32217 16167 32275 16173
rect 32217 16164 32229 16167
rect 31168 16136 32229 16164
rect 31168 16124 31174 16136
rect 32217 16133 32229 16136
rect 32263 16133 32275 16167
rect 32217 16127 32275 16133
rect 29546 15988 29552 16040
rect 29604 16028 29610 16040
rect 30009 16031 30067 16037
rect 30009 16028 30021 16031
rect 29604 16000 30021 16028
rect 29604 15988 29610 16000
rect 30009 15997 30021 16000
rect 30055 15997 30067 16031
rect 30009 15991 30067 15997
rect 30193 16031 30251 16037
rect 30193 15997 30205 16031
rect 30239 16028 30251 16031
rect 31662 16028 31668 16040
rect 30239 16000 31668 16028
rect 30239 15997 30251 16000
rect 30193 15991 30251 15997
rect 31662 15988 31668 16000
rect 31720 15988 31726 16040
rect 29549 15895 29607 15901
rect 29549 15861 29561 15895
rect 29595 15892 29607 15895
rect 30282 15892 30288 15904
rect 29595 15864 30288 15892
rect 29595 15861 29607 15864
rect 29549 15855 29607 15861
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 32493 15895 32551 15901
rect 32493 15861 32505 15895
rect 32539 15892 32551 15895
rect 77846 15892 77852 15904
rect 32539 15864 77852 15892
rect 32539 15861 32551 15864
rect 32493 15855 32551 15861
rect 77846 15852 77852 15864
rect 77904 15852 77910 15904
rect 1104 15802 78844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 78844 15802
rect 1104 15728 78844 15750
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 12492 15660 14381 15688
rect 12492 15648 12498 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 30282 15484 30288 15496
rect 30243 15456 30288 15484
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 77849 15487 77907 15493
rect 77849 15484 77861 15487
rect 64846 15456 77861 15484
rect 14274 15416 14280 15428
rect 14235 15388 14280 15416
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 30561 15351 30619 15357
rect 30561 15317 30573 15351
rect 30607 15348 30619 15351
rect 64846 15348 64874 15456
rect 77849 15453 77861 15456
rect 77895 15453 77907 15487
rect 77849 15447 77907 15453
rect 78030 15348 78036 15360
rect 30607 15320 64874 15348
rect 77991 15320 78036 15348
rect 30607 15317 30619 15320
rect 30561 15311 30619 15317
rect 78030 15308 78036 15320
rect 78088 15308 78094 15360
rect 1104 15258 78844 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 78844 15258
rect 1104 15184 78844 15206
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 14660 15076 14688 15107
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 16816 15116 16865 15144
rect 16816 15104 16822 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 18414 15144 18420 15156
rect 18375 15116 18420 15144
rect 16853 15107 16911 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 13464 15048 14688 15076
rect 13464 15017 13492 15048
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14700 14980 15209 15008
rect 14700 14968 14706 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 16298 14968 16304 15020
rect 16356 15008 16362 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16356 14980 16773 15008
rect 16356 14968 16362 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 18325 15011 18383 15017
rect 18325 15008 18337 15011
rect 17828 14980 18337 15008
rect 17828 14968 17834 14980
rect 18325 14977 18337 14980
rect 18371 14977 18383 15011
rect 18325 14971 18383 14977
rect 14182 14940 14188 14952
rect 14143 14912 14188 14940
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 14424 14912 15393 14940
rect 14424 14900 14430 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14841 14611 14875
rect 14553 14835 14611 14841
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 1452 14776 13645 14804
rect 1452 14764 1458 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 14568 14804 14596 14835
rect 15378 14804 15384 14816
rect 14568 14776 15384 14804
rect 13633 14767 13691 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 1104 14714 78844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 78844 14714
rect 1104 14640 78844 14662
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14332 14572 14657 14600
rect 14332 14560 14338 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 16298 14600 16304 14612
rect 16259 14572 16304 14600
rect 14645 14563 14703 14569
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 14461 14535 14519 14541
rect 14461 14532 14473 14535
rect 14056 14504 14473 14532
rect 14056 14492 14062 14504
rect 14461 14501 14473 14504
rect 14507 14501 14519 14535
rect 16206 14532 16212 14544
rect 16167 14504 16212 14532
rect 14461 14495 14519 14501
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 17589 14535 17647 14541
rect 17589 14501 17601 14535
rect 17635 14532 17647 14535
rect 17678 14532 17684 14544
rect 17635 14504 17684 14532
rect 17635 14501 17647 14504
rect 17589 14495 17647 14501
rect 17678 14492 17684 14504
rect 17736 14492 17742 14544
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 18371 14368 27077 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 27065 14365 27077 14368
rect 27111 14396 27123 14399
rect 77849 14399 77907 14405
rect 77849 14396 77861 14399
rect 27111 14368 35894 14396
rect 27111 14365 27123 14368
rect 27065 14359 27123 14365
rect 14182 14328 14188 14340
rect 14095 14300 14188 14328
rect 14182 14288 14188 14300
rect 14240 14328 14246 14340
rect 15841 14331 15899 14337
rect 15841 14328 15853 14331
rect 14240 14300 15853 14328
rect 14240 14288 14246 14300
rect 15841 14297 15853 14300
rect 15887 14328 15899 14331
rect 17221 14331 17279 14337
rect 17221 14328 17233 14331
rect 15887 14300 17233 14328
rect 15887 14297 15899 14300
rect 15841 14291 15899 14297
rect 17221 14297 17233 14300
rect 17267 14328 17279 14331
rect 17267 14300 18184 14328
rect 17267 14297 17279 14300
rect 17221 14291 17279 14297
rect 17681 14263 17739 14269
rect 17681 14229 17693 14263
rect 17727 14260 17739 14263
rect 17770 14260 17776 14272
rect 17727 14232 17776 14260
rect 17727 14229 17739 14232
rect 17681 14223 17739 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18156 14269 18184 14300
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 27801 14331 27859 14337
rect 27801 14328 27813 14331
rect 27304 14300 27813 14328
rect 27304 14288 27310 14300
rect 27801 14297 27813 14300
rect 27847 14297 27859 14331
rect 35866 14328 35894 14368
rect 64846 14368 77861 14396
rect 36538 14328 36544 14340
rect 35866 14300 36544 14328
rect 27801 14291 27859 14297
rect 36538 14288 36544 14300
rect 36596 14288 36602 14340
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14229 18199 14263
rect 27154 14260 27160 14272
rect 27115 14232 27160 14260
rect 18141 14223 18199 14229
rect 27154 14220 27160 14232
rect 27212 14220 27218 14272
rect 28077 14263 28135 14269
rect 28077 14229 28089 14263
rect 28123 14260 28135 14263
rect 64846 14260 64874 14368
rect 77849 14365 77861 14368
rect 77895 14365 77907 14399
rect 77849 14359 77907 14365
rect 78030 14260 78036 14272
rect 28123 14232 64874 14260
rect 77991 14232 78036 14260
rect 28123 14229 28135 14232
rect 28077 14223 28135 14229
rect 78030 14220 78036 14232
rect 78088 14220 78094 14272
rect 1104 14170 78844 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 78844 14170
rect 1104 14096 78844 14118
rect 14642 14056 14648 14068
rect 14603 14028 14648 14056
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 27157 14059 27215 14065
rect 27157 14025 27169 14059
rect 27203 14056 27215 14059
rect 27246 14056 27252 14068
rect 27203 14028 27252 14056
rect 27203 14025 27215 14028
rect 27157 14019 27215 14025
rect 27246 14016 27252 14028
rect 27304 14016 27310 14068
rect 27522 14056 27528 14068
rect 27483 14028 27528 14056
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 14182 13988 14188 14000
rect 14143 13960 14188 13988
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 26970 13948 26976 14000
rect 27028 13988 27034 14000
rect 77297 13991 77355 13997
rect 77297 13988 77309 13991
rect 27028 13960 77309 13988
rect 27028 13948 27034 13960
rect 77297 13957 77309 13960
rect 77343 13988 77355 13991
rect 77343 13960 77708 13988
rect 77343 13957 77355 13960
rect 77297 13951 77355 13957
rect 77680 13929 77708 13960
rect 77665 13923 77723 13929
rect 77665 13889 77677 13923
rect 77711 13889 77723 13923
rect 77665 13883 77723 13889
rect 27338 13812 27344 13864
rect 27396 13852 27402 13864
rect 27617 13855 27675 13861
rect 27617 13852 27629 13855
rect 27396 13824 27629 13852
rect 27396 13812 27402 13824
rect 27617 13821 27629 13824
rect 27663 13821 27675 13855
rect 27617 13815 27675 13821
rect 27709 13855 27767 13861
rect 27709 13821 27721 13855
rect 27755 13821 27767 13855
rect 27709 13815 27767 13821
rect 14458 13784 14464 13796
rect 14419 13756 14464 13784
rect 14458 13744 14464 13756
rect 14516 13744 14522 13796
rect 27154 13744 27160 13796
rect 27212 13784 27218 13796
rect 27724 13784 27752 13815
rect 27212 13756 27752 13784
rect 27212 13744 27218 13756
rect 77846 13716 77852 13728
rect 77807 13688 77852 13716
rect 77846 13676 77852 13688
rect 77904 13676 77910 13728
rect 1104 13626 78844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 78844 13626
rect 1104 13552 78844 13574
rect 26970 13512 26976 13524
rect 26931 13484 26976 13512
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 25958 13376 25964 13388
rect 25919 13348 25964 13376
rect 25958 13336 25964 13348
rect 26016 13376 26022 13388
rect 27154 13376 27160 13388
rect 26016 13348 27160 13376
rect 26016 13336 26022 13348
rect 27154 13336 27160 13348
rect 27212 13336 27218 13388
rect 25774 13308 25780 13320
rect 25735 13280 25780 13308
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 26697 13243 26755 13249
rect 26697 13240 26709 13243
rect 25424 13212 26709 13240
rect 25424 13181 25452 13212
rect 26697 13209 26709 13212
rect 26743 13209 26755 13243
rect 26697 13203 26755 13209
rect 25409 13175 25467 13181
rect 25409 13141 25421 13175
rect 25455 13141 25467 13175
rect 25409 13135 25467 13141
rect 25682 13132 25688 13184
rect 25740 13172 25746 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 25740 13144 25881 13172
rect 25740 13132 25746 13144
rect 25869 13141 25881 13144
rect 25915 13141 25927 13175
rect 25869 13135 25927 13141
rect 1104 13082 78844 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 78844 13082
rect 1104 13008 78844 13030
rect 77665 12835 77723 12841
rect 77665 12832 77677 12835
rect 77312 12804 77677 12832
rect 24762 12588 24768 12640
rect 24820 12628 24826 12640
rect 77312 12637 77340 12804
rect 77665 12801 77677 12804
rect 77711 12801 77723 12835
rect 77665 12795 77723 12801
rect 77297 12631 77355 12637
rect 77297 12628 77309 12631
rect 24820 12600 77309 12628
rect 24820 12588 24826 12600
rect 77297 12597 77309 12600
rect 77343 12597 77355 12631
rect 77846 12628 77852 12640
rect 77807 12600 77852 12628
rect 77297 12591 77355 12597
rect 77846 12588 77852 12600
rect 77904 12588 77910 12640
rect 1104 12538 78844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 78844 12538
rect 1104 12464 78844 12486
rect 24762 12424 24768 12436
rect 24723 12396 24768 12424
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 23658 12288 23664 12300
rect 23619 12260 23664 12288
rect 23658 12248 23664 12260
rect 23716 12288 23722 12300
rect 25958 12288 25964 12300
rect 23716 12260 25964 12288
rect 23716 12248 23722 12260
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 23474 12220 23480 12232
rect 23435 12192 23480 12220
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 24489 12155 24547 12161
rect 24489 12152 24501 12155
rect 23124 12124 24501 12152
rect 23124 12093 23152 12124
rect 24489 12121 24501 12124
rect 24535 12121 24547 12155
rect 24489 12115 24547 12121
rect 23109 12087 23167 12093
rect 23109 12053 23121 12087
rect 23155 12053 23167 12087
rect 23109 12047 23167 12053
rect 23569 12087 23627 12093
rect 23569 12053 23581 12087
rect 23615 12084 23627 12087
rect 24394 12084 24400 12096
rect 23615 12056 24400 12084
rect 23615 12053 23627 12056
rect 23569 12047 23627 12053
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 1104 11994 78844 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 78844 11994
rect 1104 11920 78844 11942
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21821 11883 21879 11889
rect 21821 11849 21833 11883
rect 21867 11849 21879 11883
rect 22186 11880 22192 11892
rect 22147 11852 22192 11880
rect 21821 11843 21879 11849
rect 21836 11812 21864 11843
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 23845 11815 23903 11821
rect 23845 11812 23857 11815
rect 21836 11784 23857 11812
rect 23845 11781 23857 11784
rect 23891 11781 23903 11815
rect 23845 11775 23903 11781
rect 77665 11747 77723 11753
rect 77665 11744 77677 11747
rect 64846 11716 77677 11744
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 20128 11648 20453 11676
rect 20128 11636 20134 11648
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11645 20683 11679
rect 22278 11676 22284 11688
rect 22239 11648 22284 11676
rect 20625 11639 20683 11645
rect 20640 11608 20668 11639
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 23658 11676 23664 11688
rect 22419 11648 23664 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22388 11608 22416 11639
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 20640 11580 22416 11608
rect 19978 11540 19984 11552
rect 19939 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 24121 11543 24179 11549
rect 24121 11509 24133 11543
rect 24167 11540 24179 11543
rect 64846 11540 64874 11716
rect 77665 11713 77677 11716
rect 77711 11713 77723 11747
rect 77665 11707 77723 11713
rect 77846 11608 77852 11620
rect 77807 11580 77852 11608
rect 77846 11568 77852 11580
rect 77904 11568 77910 11620
rect 24167 11512 64874 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 1104 11450 78844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 78844 11450
rect 1104 11376 78844 11398
rect 78030 11268 78036 11280
rect 77991 11240 78036 11268
rect 78030 11228 78036 11240
rect 78088 11228 78094 11280
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 23385 11135 23443 11141
rect 23385 11132 23397 11135
rect 20036 11104 23397 11132
rect 20036 11092 20042 11104
rect 23385 11101 23397 11104
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 77849 11135 77907 11141
rect 77849 11132 77861 11135
rect 23799 11104 77861 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 77849 11101 77861 11104
rect 77895 11101 77907 11135
rect 77849 11095 77907 11101
rect 1104 10906 78844 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 78844 10906
rect 1104 10832 78844 10854
rect 1104 10362 78844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 78844 10362
rect 1104 10288 78844 10310
rect 77938 10112 77944 10124
rect 77899 10084 77944 10112
rect 77938 10072 77944 10084
rect 77996 10072 78002 10124
rect 77662 10044 77668 10056
rect 77623 10016 77668 10044
rect 77662 10004 77668 10016
rect 77720 10004 77726 10056
rect 1104 9818 78844 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 78844 9818
rect 1104 9744 78844 9766
rect 1104 9274 78844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 78844 9274
rect 1104 9200 78844 9222
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 9125 9095 9183 9101
rect 9125 9092 9137 9095
rect 2924 9064 9137 9092
rect 2924 9052 2930 9064
rect 9125 9061 9137 9064
rect 9171 9061 9183 9095
rect 9125 9055 9183 9061
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 77662 8956 77668 8968
rect 77623 8928 77668 8956
rect 77662 8916 77668 8928
rect 77720 8916 77726 8968
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8386 8888 8392 8900
rect 8251 8860 8392 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 77570 8848 77576 8900
rect 77628 8888 77634 8900
rect 77941 8891 77999 8897
rect 77941 8888 77953 8891
rect 77628 8860 77953 8888
rect 77628 8848 77634 8860
rect 77941 8857 77953 8860
rect 77987 8857 77999 8891
rect 77941 8851 77999 8857
rect 1104 8730 78844 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 78844 8730
rect 1104 8656 78844 8678
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 4856 8588 8217 8616
rect 4856 8576 4862 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 8205 8579 8263 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 9030 8480 9036 8492
rect 8159 8452 9036 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9232 8452 9781 8480
rect 8754 8412 8760 8424
rect 8715 8384 8760 8412
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 9232 8421 9260 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 10502 8480 10508 8492
rect 10463 8452 10508 8480
rect 9769 8443 9827 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 9217 8415 9275 8421
rect 8864 8384 9168 8412
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 8864 8344 8892 8384
rect 6788 8316 8892 8344
rect 9033 8347 9091 8353
rect 6788 8304 6794 8316
rect 9033 8313 9045 8347
rect 9079 8313 9091 8347
rect 9140 8344 9168 8384
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 9140 8316 9965 8344
rect 9033 8307 9091 8313
rect 9953 8313 9965 8316
rect 9999 8313 10011 8347
rect 9953 8307 10011 8313
rect 9048 8276 9076 8307
rect 10042 8304 10048 8356
rect 10100 8304 10106 8356
rect 10060 8276 10088 8304
rect 9048 8248 10088 8276
rect 1104 8186 78844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 78844 8186
rect 1104 8112 78844 8134
rect 8386 8072 8392 8084
rect 8347 8044 8392 8072
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 8996 8044 9413 8072
rect 8996 8032 9002 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 10502 8072 10508 8084
rect 10367 8044 10508 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 8205 8007 8263 8013
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 9122 8004 9128 8016
rect 8251 7976 9128 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 9306 8004 9312 8016
rect 9267 7976 9312 8004
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 7973 10287 8007
rect 10229 7967 10287 7973
rect 10244 7936 10272 7967
rect 10318 7936 10324 7948
rect 10244 7908 10324 7936
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 77662 7868 77668 7880
rect 77623 7840 77668 7868
rect 77662 7828 77668 7840
rect 77720 7828 77726 7880
rect 7929 7803 7987 7809
rect 7929 7769 7941 7803
rect 7975 7800 7987 7803
rect 8754 7800 8760 7812
rect 7975 7772 8760 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 8754 7760 8760 7772
rect 8812 7800 8818 7812
rect 8941 7803 8999 7809
rect 8941 7800 8953 7803
rect 8812 7772 8953 7800
rect 8812 7760 8818 7772
rect 8941 7769 8953 7772
rect 8987 7800 8999 7803
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 8987 7772 9873 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 9861 7763 9919 7769
rect 77941 7803 77999 7809
rect 77941 7769 77953 7803
rect 77987 7800 77999 7803
rect 78030 7800 78036 7812
rect 77987 7772 78036 7800
rect 77987 7769 77999 7772
rect 77941 7763 77999 7769
rect 78030 7760 78036 7772
rect 78088 7760 78094 7812
rect 1104 7642 78844 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 78844 7642
rect 1104 7568 78844 7590
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 9088 7500 9229 7528
rect 9088 7488 9094 7500
rect 9217 7497 9229 7500
rect 9263 7497 9275 7531
rect 9217 7491 9275 7497
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 8754 7460 8760 7472
rect 8715 7432 8760 7460
rect 8754 7420 8760 7432
rect 8812 7460 8818 7472
rect 9692 7460 9720 7491
rect 8812 7432 9720 7460
rect 8812 7420 8818 7432
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 9950 7392 9956 7404
rect 9907 7364 9956 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 77202 7352 77208 7404
rect 77260 7392 77266 7404
rect 77481 7395 77539 7401
rect 77481 7392 77493 7395
rect 77260 7364 77493 7392
rect 77260 7352 77266 7364
rect 77481 7361 77493 7364
rect 77527 7361 77539 7395
rect 77481 7355 77539 7361
rect 77757 7327 77815 7333
rect 77757 7293 77769 7327
rect 77803 7324 77815 7327
rect 77846 7324 77852 7336
rect 77803 7296 77852 7324
rect 77803 7293 77815 7296
rect 77757 7287 77815 7293
rect 77846 7284 77852 7296
rect 77904 7284 77910 7336
rect 9125 7259 9183 7265
rect 9125 7225 9137 7259
rect 9171 7256 9183 7259
rect 9398 7256 9404 7268
rect 9171 7228 9404 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 9398 7216 9404 7228
rect 9456 7216 9462 7268
rect 1104 7098 78844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 78844 7098
rect 1104 7024 78844 7046
rect 1104 6554 78844 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 78844 6554
rect 1104 6480 78844 6502
rect 77478 6304 77484 6316
rect 77439 6276 77484 6304
rect 77478 6264 77484 6276
rect 77536 6264 77542 6316
rect 77386 6196 77392 6248
rect 77444 6236 77450 6248
rect 77665 6239 77723 6245
rect 77665 6236 77677 6239
rect 77444 6208 77677 6236
rect 77444 6196 77450 6208
rect 77665 6205 77677 6208
rect 77711 6205 77723 6239
rect 77665 6199 77723 6205
rect 1104 6010 78844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 78844 6010
rect 1104 5936 78844 5958
rect 1104 5466 78844 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 78844 5466
rect 1104 5392 78844 5414
rect 77478 5216 77484 5228
rect 77439 5188 77484 5216
rect 77478 5176 77484 5188
rect 77536 5176 77542 5228
rect 77665 5151 77723 5157
rect 77665 5117 77677 5151
rect 77711 5117 77723 5151
rect 77665 5111 77723 5117
rect 77478 4972 77484 5024
rect 77536 5012 77542 5024
rect 77680 5012 77708 5111
rect 77536 4984 77708 5012
rect 77536 4972 77542 4984
rect 1104 4922 78844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 78844 4922
rect 1104 4848 78844 4870
rect 77662 4604 77668 4616
rect 77623 4576 77668 4604
rect 77662 4564 77668 4576
rect 77720 4564 77726 4616
rect 77294 4496 77300 4548
rect 77352 4536 77358 4548
rect 77941 4539 77999 4545
rect 77941 4536 77953 4539
rect 77352 4508 77953 4536
rect 77352 4496 77358 4508
rect 77941 4505 77953 4508
rect 77987 4505 77999 4539
rect 77941 4499 77999 4505
rect 1104 4378 78844 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 78844 4378
rect 1104 4304 78844 4326
rect 77757 4199 77815 4205
rect 77757 4165 77769 4199
rect 77803 4196 77815 4199
rect 79042 4196 79048 4208
rect 77803 4168 79048 4196
rect 77803 4165 77815 4168
rect 77757 4159 77815 4165
rect 79042 4156 79048 4168
rect 79100 4156 79106 4208
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9582 4128 9588 4140
rect 9180 4100 9588 4128
rect 9180 4088 9186 4100
rect 9582 4088 9588 4100
rect 9640 4128 9646 4140
rect 77294 4128 77300 4140
rect 9640 4100 77300 4128
rect 9640 4088 9646 4100
rect 77294 4088 77300 4100
rect 77352 4088 77358 4140
rect 77941 4131 77999 4137
rect 77941 4097 77953 4131
rect 77987 4128 77999 4131
rect 78122 4128 78128 4140
rect 77987 4100 78128 4128
rect 77987 4097 77999 4100
rect 77941 4091 77999 4097
rect 78122 4088 78128 4100
rect 78180 4088 78186 4140
rect 1104 3834 78844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 78844 3834
rect 1104 3760 78844 3782
rect 9582 3720 9588 3732
rect 9543 3692 9588 3720
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9600 3584 9628 3680
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 21358 3652 21364 3664
rect 14056 3624 21364 3652
rect 14056 3612 14062 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 9140 3556 9628 3584
rect 9140 3525 9168 3556
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 77754 3584 77760 3596
rect 9732 3556 77760 3584
rect 9732 3544 9738 3556
rect 77754 3544 77760 3556
rect 77812 3544 77818 3596
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8435 3488 8953 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9950 3516 9956 3528
rect 9355 3488 9812 3516
rect 9911 3488 9956 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9784 3389 9812 3488
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3516 16543 3519
rect 16666 3516 16672 3528
rect 16531 3488 16672 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 9968 3448 9996 3476
rect 15856 3448 15884 3479
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 50982 3516 50988 3528
rect 20824 3488 50988 3516
rect 20824 3448 20852 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 77662 3516 77668 3528
rect 77623 3488 77668 3516
rect 77662 3476 77668 3488
rect 77720 3476 77726 3528
rect 9968 3420 20852 3448
rect 21358 3408 21364 3460
rect 21416 3448 21422 3460
rect 77386 3448 77392 3460
rect 21416 3420 77392 3448
rect 21416 3408 21422 3420
rect 77386 3408 77392 3420
rect 77444 3408 77450 3460
rect 77938 3448 77944 3460
rect 77899 3420 77944 3448
rect 77938 3408 77944 3420
rect 77996 3408 78002 3460
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 8168 3352 8217 3380
rect 8168 3340 8174 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 8205 3343 8263 3349
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 9858 3380 9864 3392
rect 9815 3352 9864 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14277 3383 14335 3389
rect 14277 3380 14289 3383
rect 13872 3352 14289 3380
rect 13872 3340 13878 3352
rect 14277 3349 14289 3352
rect 14323 3349 14335 3383
rect 14277 3343 14335 3349
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 15657 3383 15715 3389
rect 15657 3380 15669 3383
rect 15160 3352 15669 3380
rect 15160 3340 15166 3352
rect 15657 3349 15669 3352
rect 15703 3349 15715 3383
rect 15657 3343 15715 3349
rect 16301 3383 16359 3389
rect 16301 3349 16313 3383
rect 16347 3380 16359 3383
rect 16574 3380 16580 3392
rect 16347 3352 16580 3380
rect 16347 3349 16359 3352
rect 16301 3343 16359 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 76282 3340 76288 3392
rect 76340 3380 76346 3392
rect 78030 3380 78036 3392
rect 76340 3352 78036 3380
rect 76340 3340 76346 3352
rect 78030 3340 78036 3352
rect 78088 3340 78094 3392
rect 1104 3290 78844 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 78844 3290
rect 1104 3216 78844 3238
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 16206 3176 16212 3188
rect 16167 3148 16212 3176
rect 16206 3136 16212 3148
rect 16264 3176 16270 3188
rect 16666 3176 16672 3188
rect 16264 3148 16574 3176
rect 16627 3148 16672 3176
rect 16264 3136 16270 3148
rect 9309 3111 9367 3117
rect 9309 3108 9321 3111
rect 8404 3080 9321 3108
rect 8404 3049 8432 3080
rect 9309 3077 9321 3080
rect 9355 3077 9367 3111
rect 14016 3108 14044 3136
rect 14016 3080 14596 3108
rect 9309 3071 9367 3077
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 9122 3040 9128 3052
rect 9083 3012 9128 3040
rect 8389 3003 8447 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 10042 3040 10048 3052
rect 9955 3012 10048 3040
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10275 3012 10701 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14274 3040 14280 3052
rect 13771 3012 14280 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14568 3049 14596 3080
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14700 3012 14749 3040
rect 14700 3000 14706 3012
rect 14737 3009 14749 3012
rect 14783 3040 14795 3043
rect 15102 3040 15108 3052
rect 14783 3012 15108 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 15102 3000 15108 3012
rect 15160 3040 15166 3052
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15160 3012 15301 3040
rect 15160 3000 15166 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 8987 2944 9413 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 9401 2941 9413 2944
rect 9447 2972 9459 2975
rect 9858 2972 9864 2984
rect 9447 2944 9864 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 10060 2972 10088 3000
rect 15304 2972 15332 3003
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 16546 3040 16574 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 76282 3176 76288 3188
rect 16868 3148 76288 3176
rect 16868 3049 16896 3148
rect 76282 3136 76288 3148
rect 76340 3136 76346 3188
rect 76926 3176 76932 3188
rect 76887 3148 76932 3176
rect 76926 3136 76932 3148
rect 76984 3136 76990 3188
rect 77938 3108 77944 3120
rect 17604 3080 77944 3108
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 15436 3012 15481 3040
rect 16546 3012 16865 3040
rect 15436 3000 15442 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 10060 2944 15240 2972
rect 15304 2944 17049 2972
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 10505 2907 10563 2913
rect 10505 2904 10517 2907
rect 7616 2876 10517 2904
rect 7616 2864 7622 2876
rect 10505 2873 10517 2876
rect 10551 2873 10563 2907
rect 10505 2867 10563 2873
rect 13541 2907 13599 2913
rect 13541 2873 13553 2907
rect 13587 2904 13599 2907
rect 15102 2904 15108 2916
rect 13587 2876 15108 2904
rect 13587 2873 13599 2876
rect 13541 2867 13599 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 15212 2904 15240 2944
rect 17037 2941 17049 2944
rect 17083 2972 17095 2975
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17083 2944 17509 2972
rect 17083 2941 17095 2944
rect 17037 2935 17095 2941
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 17604 2904 17632 3080
rect 77938 3068 77944 3080
rect 77996 3068 78002 3120
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17865 3043 17923 3049
rect 17736 3012 17829 3040
rect 17736 3000 17742 3012
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 17911 3012 18521 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 41325 3043 41383 3049
rect 41325 3009 41337 3043
rect 41371 3040 41383 3043
rect 41506 3040 41512 3052
rect 41371 3012 41512 3040
rect 41371 3009 41383 3012
rect 41325 3003 41383 3009
rect 41506 3000 41512 3012
rect 41564 3000 41570 3052
rect 76837 3043 76895 3049
rect 76837 3009 76849 3043
rect 76883 3040 76895 3043
rect 77110 3040 77116 3052
rect 76883 3012 77116 3040
rect 76883 3009 76895 3012
rect 76837 3003 76895 3009
rect 77110 3000 77116 3012
rect 77168 3000 77174 3052
rect 77481 3043 77539 3049
rect 77481 3009 77493 3043
rect 77527 3009 77539 3043
rect 77754 3040 77760 3052
rect 77715 3012 77760 3040
rect 77481 3003 77539 3009
rect 17696 2972 17724 3000
rect 17696 2944 18276 2972
rect 18248 2913 18276 2944
rect 40954 2932 40960 2984
rect 41012 2972 41018 2984
rect 41049 2975 41107 2981
rect 41049 2972 41061 2975
rect 41012 2944 41061 2972
rect 41012 2932 41018 2944
rect 41049 2941 41061 2944
rect 41095 2941 41107 2975
rect 41049 2935 41107 2941
rect 77018 2932 77024 2984
rect 77076 2972 77082 2984
rect 77496 2972 77524 3003
rect 77754 3000 77760 3012
rect 77812 3000 77818 3052
rect 77076 2944 77524 2972
rect 77076 2932 77082 2944
rect 15212 2876 17632 2904
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2904 18291 2907
rect 77570 2904 77576 2916
rect 18279 2876 77576 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 77570 2864 77576 2876
rect 77628 2864 77634 2916
rect 8202 2836 8208 2848
rect 8163 2808 8208 2836
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 8444 2808 9781 2836
rect 8444 2796 8450 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 15565 2839 15623 2845
rect 15565 2836 15577 2839
rect 14148 2808 15577 2836
rect 14148 2796 14154 2808
rect 15565 2805 15577 2808
rect 15611 2805 15623 2839
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 15565 2799 15623 2805
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 1104 2746 78844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 78844 2746
rect 1104 2672 78844 2694
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 1412 2604 13369 2632
rect 1412 2437 1440 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 13357 2595 13415 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 20070 2632 20076 2644
rect 20031 2604 20076 2632
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 21913 2635 21971 2641
rect 21913 2601 21925 2635
rect 21959 2632 21971 2635
rect 22278 2632 22284 2644
rect 21959 2604 22284 2632
rect 21959 2601 21971 2604
rect 21913 2595 21971 2601
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 24394 2632 24400 2644
rect 24355 2604 24400 2632
rect 24394 2592 24400 2604
rect 24452 2592 24458 2644
rect 25682 2592 25688 2644
rect 25740 2632 25746 2644
rect 25777 2635 25835 2641
rect 25777 2632 25789 2635
rect 25740 2604 25789 2632
rect 25740 2592 25746 2604
rect 25777 2601 25789 2604
rect 25823 2601 25835 2635
rect 25777 2595 25835 2601
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 27709 2635 27767 2641
rect 27709 2632 27721 2635
rect 27396 2604 27721 2632
rect 27396 2592 27402 2604
rect 27709 2601 27721 2604
rect 27755 2601 27767 2635
rect 29546 2632 29552 2644
rect 29507 2604 29552 2632
rect 27709 2595 27767 2601
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 31570 2592 31576 2644
rect 31628 2632 31634 2644
rect 32125 2635 32183 2641
rect 32125 2632 32137 2635
rect 31628 2604 32137 2632
rect 31628 2592 31634 2604
rect 32125 2601 32137 2604
rect 32171 2601 32183 2635
rect 32125 2595 32183 2601
rect 46658 2592 46664 2644
rect 46716 2632 46722 2644
rect 47811 2635 47869 2641
rect 47811 2632 47823 2635
rect 46716 2604 47823 2632
rect 46716 2592 46722 2604
rect 47811 2601 47823 2604
rect 47857 2601 47869 2635
rect 47811 2595 47869 2601
rect 49053 2635 49111 2641
rect 49053 2601 49065 2635
rect 49099 2632 49111 2635
rect 49142 2632 49148 2644
rect 49099 2604 49148 2632
rect 49099 2601 49111 2604
rect 49053 2595 49111 2601
rect 49142 2592 49148 2604
rect 49200 2592 49206 2644
rect 50706 2632 50712 2644
rect 50667 2604 50712 2632
rect 50706 2592 50712 2604
rect 50764 2592 50770 2644
rect 52914 2632 52920 2644
rect 52875 2604 52920 2632
rect 52914 2592 52920 2604
rect 52972 2592 52978 2644
rect 54570 2632 54576 2644
rect 54531 2604 54576 2632
rect 54570 2592 54576 2604
rect 54628 2592 54634 2644
rect 56410 2632 56416 2644
rect 56371 2604 56416 2632
rect 56410 2592 56416 2604
rect 56468 2592 56474 2644
rect 58342 2632 58348 2644
rect 58303 2604 58348 2632
rect 58342 2592 58348 2604
rect 58400 2592 58406 2644
rect 61838 2592 61844 2644
rect 61896 2632 61902 2644
rect 62117 2635 62175 2641
rect 62117 2632 62129 2635
rect 61896 2604 62129 2632
rect 61896 2592 61902 2604
rect 62117 2601 62129 2604
rect 62163 2601 62175 2635
rect 62117 2595 62175 2601
rect 64049 2635 64107 2641
rect 64049 2601 64061 2635
rect 64095 2632 64107 2635
rect 64138 2632 64144 2644
rect 64095 2604 64144 2632
rect 64095 2601 64107 2604
rect 64049 2595 64107 2601
rect 64138 2592 64144 2604
rect 64196 2592 64202 2644
rect 65981 2635 66039 2641
rect 65981 2601 65993 2635
rect 66027 2632 66039 2635
rect 66070 2632 66076 2644
rect 66027 2604 66076 2632
rect 66027 2601 66039 2604
rect 65981 2595 66039 2601
rect 66070 2592 66076 2604
rect 66128 2592 66134 2644
rect 68370 2632 68376 2644
rect 68331 2604 68376 2632
rect 68370 2592 68376 2604
rect 68428 2592 68434 2644
rect 69753 2635 69811 2641
rect 69753 2601 69765 2635
rect 69799 2632 69811 2635
rect 69842 2632 69848 2644
rect 69799 2604 69848 2632
rect 69799 2601 69811 2604
rect 69753 2595 69811 2601
rect 69842 2592 69848 2604
rect 69900 2592 69906 2644
rect 71406 2592 71412 2644
rect 71464 2632 71470 2644
rect 71685 2635 71743 2641
rect 71685 2632 71697 2635
rect 71464 2604 71697 2632
rect 71464 2592 71470 2604
rect 71685 2601 71697 2604
rect 71731 2601 71743 2635
rect 73614 2632 73620 2644
rect 73575 2604 73620 2632
rect 71685 2595 71743 2601
rect 73614 2592 73620 2604
rect 73672 2592 73678 2644
rect 75178 2592 75184 2644
rect 75236 2632 75242 2644
rect 75273 2635 75331 2641
rect 75273 2632 75285 2635
rect 75236 2604 75285 2632
rect 75236 2592 75242 2604
rect 75273 2601 75285 2604
rect 75319 2601 75331 2635
rect 75273 2595 75331 2601
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 6886 2536 7481 2564
rect 6886 2496 6914 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 77846 2564 77852 2576
rect 7469 2527 7527 2533
rect 14936 2536 77852 2564
rect 8386 2496 8392 2508
rect 4816 2468 6914 2496
rect 7668 2468 8392 2496
rect 4816 2437 4844 2468
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7558 2428 7564 2440
rect 6779 2400 7564 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 2884 2360 2912 2391
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7668 2437 7696 2468
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2496 9551 2499
rect 10137 2499 10195 2505
rect 9539 2468 9996 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 9968 2440 9996 2468
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 13814 2496 13820 2508
rect 10183 2468 11744 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 7653 2391 7711 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10318 2428 10324 2440
rect 10008 2400 10324 2428
rect 10008 2388 10014 2400
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11716 2437 11744 2468
rect 12452 2468 13820 2496
rect 12452 2437 12480 2468
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 14642 2496 14648 2508
rect 14603 2468 14648 2496
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 11701 2431 11759 2437
rect 10643 2400 11560 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 8202 2360 8208 2372
rect 2884 2332 8208 2360
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 992 2264 1593 2292
rect 992 2252 998 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 2832 2264 3065 2292
rect 2832 2252 2838 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 4764 2264 4997 2292
rect 4764 2252 4770 2264
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6696 2264 6929 2292
rect 6696 2252 6702 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 6917 2255 6975 2261
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8478 2292 8484 2304
rect 8343 2264 8484 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 11532 2301 11560 2400
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 14090 2428 14096 2440
rect 13587 2400 14096 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 14458 2388 14464 2400
rect 14516 2428 14522 2440
rect 14936 2437 14964 2536
rect 77846 2524 77852 2536
rect 77904 2524 77910 2576
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 76745 2499 76803 2505
rect 76745 2496 76757 2499
rect 15436 2468 76757 2496
rect 15436 2456 15442 2468
rect 76745 2465 76757 2468
rect 76791 2465 76803 2499
rect 76745 2459 76803 2465
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14516 2400 14933 2428
rect 14516 2388 14522 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 15102 2428 15108 2440
rect 15063 2400 15108 2428
rect 14921 2391 14979 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16632 2400 16681 2428
rect 16632 2388 16638 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18322 2428 18328 2440
rect 18187 2400 18328 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21876 2400 22109 2428
rect 21876 2388 21882 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23808 2400 24593 2428
rect 23808 2388 23814 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25740 2400 25973 2428
rect 25740 2388 25746 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 27893 2431 27951 2437
rect 27893 2428 27905 2431
rect 27672 2400 27905 2428
rect 27672 2388 27678 2400
rect 27893 2397 27905 2400
rect 27939 2397 27951 2431
rect 27893 2391 27951 2397
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29512 2400 29745 2428
rect 29512 2388 29518 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31444 2400 32321 2428
rect 31444 2388 31450 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 33318 2428 33324 2440
rect 33279 2400 33324 2428
rect 32309 2391 32367 2397
rect 33318 2388 33324 2400
rect 33376 2388 33382 2440
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 35158 2388 35164 2440
rect 35216 2428 35222 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35216 2400 35265 2428
rect 35216 2388 35222 2400
rect 35253 2397 35265 2400
rect 35299 2397 35311 2431
rect 35526 2428 35532 2440
rect 35487 2400 35532 2428
rect 35253 2391 35311 2397
rect 35526 2388 35532 2400
rect 35584 2388 35590 2440
rect 37090 2388 37096 2440
rect 37148 2428 37154 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 37148 2400 37289 2428
rect 37148 2388 37154 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37550 2428 37556 2440
rect 37511 2400 37556 2428
rect 37277 2391 37335 2397
rect 37550 2388 37556 2400
rect 37608 2388 37614 2440
rect 39022 2388 39028 2440
rect 39080 2428 39086 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39080 2400 39865 2428
rect 39080 2388 39086 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 40126 2428 40132 2440
rect 40087 2400 40132 2428
rect 39853 2391 39911 2397
rect 40126 2388 40132 2400
rect 40184 2388 40190 2440
rect 42794 2388 42800 2440
rect 42852 2428 42858 2440
rect 42889 2431 42947 2437
rect 42889 2428 42901 2431
rect 42852 2400 42901 2428
rect 42852 2388 42858 2400
rect 42889 2397 42901 2400
rect 42935 2397 42947 2431
rect 43162 2428 43168 2440
rect 43123 2400 43168 2428
rect 42889 2391 42947 2397
rect 43162 2388 43168 2400
rect 43220 2388 43226 2440
rect 44726 2388 44732 2440
rect 44784 2428 44790 2440
rect 45005 2431 45063 2437
rect 45005 2428 45017 2431
rect 44784 2400 45017 2428
rect 44784 2388 44790 2400
rect 45005 2397 45017 2400
rect 45051 2397 45063 2431
rect 45278 2428 45284 2440
rect 45239 2400 45284 2428
rect 45005 2391 45063 2397
rect 45278 2388 45284 2400
rect 45336 2388 45342 2440
rect 46658 2388 46664 2440
rect 46716 2428 46722 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 46716 2400 47593 2428
rect 46716 2388 46722 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 60734 2428 60740 2440
rect 60695 2400 60740 2428
rect 47581 2391 47639 2397
rect 60734 2388 60740 2400
rect 60792 2388 60798 2440
rect 73338 2388 73344 2440
rect 73396 2428 73402 2440
rect 73433 2431 73491 2437
rect 73433 2428 73445 2431
rect 73396 2400 73445 2428
rect 73396 2388 73402 2400
rect 73433 2397 73445 2400
rect 73479 2397 73491 2431
rect 73433 2391 73491 2397
rect 75089 2431 75147 2437
rect 75089 2397 75101 2431
rect 75135 2428 75147 2431
rect 75178 2428 75184 2440
rect 75135 2400 75184 2428
rect 75135 2397 75147 2400
rect 75089 2391 75147 2397
rect 75178 2388 75184 2400
rect 75236 2388 75242 2440
rect 76558 2428 76564 2440
rect 76519 2400 76564 2428
rect 76558 2388 76564 2400
rect 76616 2388 76622 2440
rect 77202 2388 77208 2440
rect 77260 2428 77266 2440
rect 77481 2431 77539 2437
rect 77481 2428 77493 2431
rect 77260 2400 77493 2428
rect 77260 2388 77266 2400
rect 77481 2397 77493 2400
rect 77527 2397 77539 2431
rect 77481 2391 77539 2397
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 14332 2332 15332 2360
rect 14332 2320 14338 2332
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10468 2264 10793 2292
rect 10468 2252 10474 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 11517 2295 11575 2301
rect 11517 2261 11529 2295
rect 11563 2261 11575 2295
rect 11517 2255 11575 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 15304 2301 15332 2332
rect 48498 2320 48504 2372
rect 48556 2360 48562 2372
rect 48961 2363 49019 2369
rect 48961 2360 48973 2363
rect 48556 2332 48973 2360
rect 48556 2320 48562 2332
rect 48961 2329 48973 2332
rect 49007 2329 49019 2363
rect 50614 2360 50620 2372
rect 50575 2332 50620 2360
rect 48961 2323 49019 2329
rect 50614 2320 50620 2332
rect 50672 2320 50678 2372
rect 52362 2320 52368 2372
rect 52420 2360 52426 2372
rect 52825 2363 52883 2369
rect 52825 2360 52837 2363
rect 52420 2332 52837 2360
rect 52420 2320 52426 2332
rect 52825 2329 52837 2332
rect 52871 2329 52883 2363
rect 52825 2323 52883 2329
rect 54294 2320 54300 2372
rect 54352 2360 54358 2372
rect 54481 2363 54539 2369
rect 54481 2360 54493 2363
rect 54352 2332 54493 2360
rect 54352 2320 54358 2332
rect 54481 2329 54493 2332
rect 54527 2329 54539 2363
rect 54481 2323 54539 2329
rect 56134 2320 56140 2372
rect 56192 2360 56198 2372
rect 56321 2363 56379 2369
rect 56321 2360 56333 2363
rect 56192 2332 56333 2360
rect 56192 2320 56198 2332
rect 56321 2329 56333 2332
rect 56367 2329 56379 2363
rect 56321 2323 56379 2329
rect 58066 2320 58072 2372
rect 58124 2360 58130 2372
rect 58253 2363 58311 2369
rect 58253 2360 58265 2363
rect 58124 2332 58265 2360
rect 58124 2320 58130 2332
rect 58253 2329 58265 2332
rect 58299 2329 58311 2363
rect 58253 2323 58311 2329
rect 59998 2320 60004 2372
rect 60056 2360 60062 2372
rect 60553 2363 60611 2369
rect 60553 2360 60565 2363
rect 60056 2332 60565 2360
rect 60056 2320 60062 2332
rect 60553 2329 60565 2332
rect 60599 2329 60611 2363
rect 60553 2323 60611 2329
rect 61838 2320 61844 2372
rect 61896 2360 61902 2372
rect 62025 2363 62083 2369
rect 62025 2360 62037 2363
rect 61896 2332 62037 2360
rect 61896 2320 61902 2332
rect 62025 2329 62037 2332
rect 62071 2329 62083 2363
rect 62025 2323 62083 2329
rect 63770 2320 63776 2372
rect 63828 2360 63834 2372
rect 63957 2363 64015 2369
rect 63957 2360 63969 2363
rect 63828 2332 63969 2360
rect 63828 2320 63834 2332
rect 63957 2329 63969 2332
rect 64003 2329 64015 2363
rect 63957 2323 64015 2329
rect 65702 2320 65708 2372
rect 65760 2360 65766 2372
rect 65889 2363 65947 2369
rect 65889 2360 65901 2363
rect 65760 2332 65901 2360
rect 65760 2320 65766 2332
rect 65889 2329 65901 2332
rect 65935 2329 65947 2363
rect 65889 2323 65947 2329
rect 67634 2320 67640 2372
rect 67692 2360 67698 2372
rect 68281 2363 68339 2369
rect 68281 2360 68293 2363
rect 67692 2332 68293 2360
rect 67692 2320 67698 2332
rect 68281 2329 68293 2332
rect 68327 2329 68339 2363
rect 68281 2323 68339 2329
rect 69474 2320 69480 2372
rect 69532 2360 69538 2372
rect 69661 2363 69719 2369
rect 69661 2360 69673 2363
rect 69532 2332 69673 2360
rect 69532 2320 69538 2332
rect 69661 2329 69673 2332
rect 69707 2329 69719 2363
rect 69661 2323 69719 2329
rect 71406 2320 71412 2372
rect 71464 2360 71470 2372
rect 71593 2363 71651 2369
rect 71593 2360 71605 2363
rect 71464 2332 71605 2360
rect 71464 2320 71470 2332
rect 71593 2329 71605 2332
rect 71639 2329 71651 2363
rect 77754 2360 77760 2372
rect 77715 2332 77760 2360
rect 71593 2323 71651 2329
rect 77754 2320 77760 2332
rect 77812 2320 77818 2372
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 12400 2264 12633 2292
rect 12400 2252 12406 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16172 2264 16865 2292
rect 16172 2252 16178 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 1104 2202 78844 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 78844 2202
rect 1104 2128 78844 2150
rect 9950 1980 9956 2032
rect 10008 2020 10014 2032
rect 77478 2020 77484 2032
rect 10008 1992 77484 2020
rect 10008 1980 10014 1992
rect 77478 1980 77484 1992
rect 77536 1980 77542 2032
rect 9122 1912 9128 1964
rect 9180 1952 9186 1964
rect 77754 1952 77760 1964
rect 9180 1924 77760 1952
rect 9180 1912 9186 1924
rect 77754 1912 77760 1924
rect 77812 1912 77818 1964
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 77208 37408 77260 37460
rect 77852 37451 77904 37460
rect 77852 37417 77861 37451
rect 77861 37417 77895 37451
rect 77895 37417 77904 37451
rect 77852 37408 77904 37417
rect 20352 37315 20404 37324
rect 20352 37281 20361 37315
rect 20361 37281 20395 37315
rect 20395 37281 20404 37315
rect 20352 37272 20404 37281
rect 22192 37315 22244 37324
rect 22192 37281 22201 37315
rect 22201 37281 22235 37315
rect 22235 37281 22244 37315
rect 22192 37272 22244 37281
rect 23480 37272 23532 37324
rect 25780 37272 25832 37324
rect 27528 37272 27580 37324
rect 29460 37272 29512 37324
rect 31392 37272 31444 37324
rect 35348 37272 35400 37324
rect 37096 37272 37148 37324
rect 39028 37272 39080 37324
rect 42800 37272 42852 37324
rect 44732 37272 44784 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 2872 37247 2924 37256
rect 2872 37213 2881 37247
rect 2881 37213 2915 37247
rect 2915 37213 2924 37247
rect 2872 37204 2924 37213
rect 4804 37247 4856 37256
rect 4804 37213 4813 37247
rect 4813 37213 4847 37247
rect 4847 37213 4856 37247
rect 4804 37204 4856 37213
rect 6736 37247 6788 37256
rect 6736 37213 6745 37247
rect 6745 37213 6779 37247
rect 6779 37213 6788 37247
rect 6736 37204 6788 37213
rect 8300 37204 8352 37256
rect 10600 37204 10652 37256
rect 12440 37247 12492 37256
rect 12440 37213 12449 37247
rect 12449 37213 12483 37247
rect 12483 37213 12492 37247
rect 12440 37204 12492 37213
rect 14372 37247 14424 37256
rect 14372 37213 14381 37247
rect 14381 37213 14415 37247
rect 14415 37213 14424 37247
rect 14372 37204 14424 37213
rect 16764 37204 16816 37256
rect 18420 37204 18472 37256
rect 19984 37204 20036 37256
rect 21824 37204 21876 37256
rect 23756 37204 23808 37256
rect 25688 37204 25740 37256
rect 27620 37204 27672 37256
rect 29920 37204 29972 37256
rect 32404 37247 32456 37256
rect 32404 37213 32413 37247
rect 32413 37213 32447 37247
rect 32447 37213 32456 37247
rect 32404 37204 32456 37213
rect 35440 37204 35492 37256
rect 37648 37204 37700 37256
rect 40224 37204 40276 37256
rect 44824 37204 44876 37256
rect 46664 37204 46716 37256
rect 48504 37204 48556 37256
rect 50436 37204 50488 37256
rect 52460 37204 52512 37256
rect 54300 37204 54352 37256
rect 56140 37204 56192 37256
rect 58072 37204 58124 37256
rect 60004 37204 60056 37256
rect 61844 37204 61896 37256
rect 63776 37204 63828 37256
rect 65984 37247 66036 37256
rect 65984 37213 65993 37247
rect 65993 37213 66027 37247
rect 66027 37213 66036 37247
rect 65984 37204 66036 37213
rect 67640 37204 67692 37256
rect 69480 37204 69532 37256
rect 71412 37204 71464 37256
rect 73344 37204 73396 37256
rect 75184 37204 75236 37256
rect 42800 37136 42852 37188
rect 74724 37136 74776 37188
rect 76932 37247 76984 37256
rect 76932 37213 76941 37247
rect 76941 37213 76975 37247
rect 76975 37213 76984 37247
rect 76932 37204 76984 37213
rect 940 37068 992 37120
rect 2780 37068 2832 37120
rect 4712 37068 4764 37120
rect 6644 37068 6696 37120
rect 8484 37068 8536 37120
rect 10416 37068 10468 37120
rect 12348 37068 12400 37120
rect 14280 37068 14332 37120
rect 16580 37068 16632 37120
rect 18052 37068 18104 37120
rect 46572 37068 46624 37120
rect 48872 37068 48924 37120
rect 50804 37068 50856 37120
rect 52460 37068 52512 37120
rect 54392 37111 54444 37120
rect 54392 37077 54401 37111
rect 54401 37077 54435 37111
rect 54435 37077 54444 37111
rect 54392 37068 54444 37077
rect 56048 37068 56100 37120
rect 58440 37068 58492 37120
rect 60648 37068 60700 37120
rect 61936 37111 61988 37120
rect 61936 37077 61945 37111
rect 61945 37077 61979 37111
rect 61979 37077 61988 37111
rect 61936 37068 61988 37077
rect 63868 37111 63920 37120
rect 63868 37077 63877 37111
rect 63877 37077 63911 37111
rect 63911 37077 63920 37111
rect 63868 37068 63920 37077
rect 66168 37068 66220 37120
rect 68192 37111 68244 37120
rect 68192 37077 68201 37111
rect 68201 37077 68235 37111
rect 68235 37077 68244 37111
rect 68192 37068 68244 37077
rect 69572 37111 69624 37120
rect 69572 37077 69581 37111
rect 69581 37077 69615 37111
rect 69615 37077 69624 37111
rect 69572 37068 69624 37077
rect 71504 37111 71556 37120
rect 71504 37077 71513 37111
rect 71513 37077 71547 37111
rect 71547 37077 71556 37111
rect 71504 37068 71556 37077
rect 73712 37068 73764 37120
rect 75092 37068 75144 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 73712 36907 73764 36916
rect 73712 36873 73721 36907
rect 73721 36873 73755 36907
rect 73755 36873 73764 36907
rect 73712 36864 73764 36873
rect 74724 36907 74776 36916
rect 74724 36873 74733 36907
rect 74733 36873 74767 36907
rect 74767 36873 74776 36907
rect 74724 36864 74776 36873
rect 75092 36907 75144 36916
rect 75092 36873 75101 36907
rect 75101 36873 75135 36907
rect 75135 36873 75144 36907
rect 75092 36864 75144 36873
rect 76748 36864 76800 36916
rect 33324 36728 33376 36780
rect 40960 36728 41012 36780
rect 76196 36728 76248 36780
rect 77668 36771 77720 36780
rect 77668 36737 77677 36771
rect 77677 36737 77711 36771
rect 77711 36737 77720 36771
rect 77668 36728 77720 36737
rect 41328 36703 41380 36712
rect 41328 36669 41337 36703
rect 41337 36669 41371 36703
rect 41371 36669 41380 36703
rect 41328 36660 41380 36669
rect 73620 36660 73672 36712
rect 73988 36703 74040 36712
rect 73988 36669 73997 36703
rect 73997 36669 74031 36703
rect 74031 36669 74040 36703
rect 75184 36703 75236 36712
rect 73988 36660 74040 36669
rect 33324 36592 33376 36644
rect 75184 36669 75193 36703
rect 75193 36669 75227 36703
rect 75227 36669 75236 36703
rect 75184 36660 75236 36669
rect 77852 36635 77904 36644
rect 77852 36601 77861 36635
rect 77861 36601 77895 36635
rect 77895 36601 77904 36635
rect 77852 36592 77904 36601
rect 73804 36524 73856 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 77668 36184 77720 36236
rect 73804 36159 73856 36168
rect 73804 36125 73813 36159
rect 73813 36125 73847 36159
rect 73847 36125 73856 36159
rect 73804 36116 73856 36125
rect 77116 36116 77168 36168
rect 73160 36048 73212 36100
rect 76748 35980 76800 36032
rect 78036 36023 78088 36032
rect 78036 35989 78045 36023
rect 78045 35989 78079 36023
rect 78079 35989 78088 36023
rect 78036 35980 78088 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 71504 35819 71556 35828
rect 71504 35785 71513 35819
rect 71513 35785 71547 35819
rect 71547 35785 71556 35819
rect 71504 35776 71556 35785
rect 73160 35776 73212 35828
rect 71412 35572 71464 35624
rect 73252 35708 73304 35760
rect 73988 35708 74040 35760
rect 79048 35640 79100 35692
rect 77760 35479 77812 35488
rect 77760 35445 77769 35479
rect 77769 35445 77803 35479
rect 77803 35445 77812 35479
rect 77760 35436 77812 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 77852 35071 77904 35080
rect 77852 35037 77861 35071
rect 77861 35037 77895 35071
rect 77895 35037 77904 35071
rect 77852 35028 77904 35037
rect 78036 34935 78088 34944
rect 78036 34901 78045 34935
rect 78045 34901 78079 34935
rect 78079 34901 78088 34935
rect 78036 34892 78088 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 69572 34731 69624 34740
rect 69572 34697 69581 34731
rect 69581 34697 69615 34731
rect 69615 34697 69624 34731
rect 69572 34688 69624 34697
rect 76932 34688 76984 34740
rect 69848 34552 69900 34604
rect 77852 34620 77904 34672
rect 77208 34595 77260 34604
rect 77208 34561 77217 34595
rect 77217 34561 77251 34595
rect 77251 34561 77260 34595
rect 77208 34552 77260 34561
rect 77300 34552 77352 34604
rect 68376 34416 68428 34468
rect 73252 34416 73304 34468
rect 77852 34391 77904 34400
rect 77852 34357 77861 34391
rect 77861 34357 77895 34391
rect 77895 34357 77904 34391
rect 77852 34348 77904 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 76196 34187 76248 34196
rect 76196 34153 76205 34187
rect 76205 34153 76239 34187
rect 76239 34153 76248 34187
rect 76196 34144 76248 34153
rect 77208 34144 77260 34196
rect 68376 34051 68428 34060
rect 68376 34017 68385 34051
rect 68385 34017 68419 34051
rect 68419 34017 68428 34051
rect 68376 34008 68428 34017
rect 77116 34008 77168 34060
rect 68192 33940 68244 33992
rect 77208 33940 77260 33992
rect 76932 33872 76984 33924
rect 67732 33847 67784 33856
rect 67732 33813 67741 33847
rect 67741 33813 67775 33847
rect 67775 33813 67784 33847
rect 67732 33804 67784 33813
rect 68376 33804 68428 33856
rect 76748 33804 76800 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 73252 33600 73304 33652
rect 77208 33643 77260 33652
rect 77208 33609 77217 33643
rect 77217 33609 77251 33643
rect 77251 33609 77260 33643
rect 77208 33600 77260 33609
rect 77760 33600 77812 33652
rect 67732 33464 67784 33516
rect 68928 33464 68980 33516
rect 77944 33532 77996 33584
rect 78128 33464 78180 33516
rect 77300 33396 77352 33448
rect 77116 33328 77168 33380
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 78036 33031 78088 33040
rect 78036 32997 78045 33031
rect 78045 32997 78079 33031
rect 78079 32997 78088 33031
rect 78036 32988 78088 32997
rect 76196 32852 76248 32904
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 65984 32419 66036 32428
rect 65984 32385 65993 32419
rect 65993 32385 66027 32419
rect 66027 32385 66036 32419
rect 65984 32376 66036 32385
rect 77668 32419 77720 32428
rect 77668 32385 77677 32419
rect 77677 32385 77711 32419
rect 77711 32385 77720 32419
rect 77668 32376 77720 32385
rect 76196 32172 76248 32224
rect 77852 32215 77904 32224
rect 77852 32181 77861 32215
rect 77861 32181 77895 32215
rect 77895 32181 77904 32215
rect 77852 32172 77904 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 65984 31968 66036 32020
rect 49976 31764 50028 31816
rect 68928 31900 68980 31952
rect 63040 31807 63092 31816
rect 63040 31773 63049 31807
rect 63049 31773 63083 31807
rect 63083 31773 63092 31807
rect 63040 31764 63092 31773
rect 63500 31764 63552 31816
rect 77668 31764 77720 31816
rect 66168 31696 66220 31748
rect 66076 31671 66128 31680
rect 66076 31637 66085 31671
rect 66085 31637 66119 31671
rect 66119 31637 66128 31671
rect 66076 31628 66128 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 61936 31467 61988 31476
rect 61936 31433 61945 31467
rect 61945 31433 61979 31467
rect 61979 31433 61988 31467
rect 61936 31424 61988 31433
rect 63500 31467 63552 31476
rect 63500 31433 63509 31467
rect 63509 31433 63543 31467
rect 63543 31433 63552 31467
rect 63500 31424 63552 31433
rect 63868 31467 63920 31476
rect 63868 31433 63877 31467
rect 63877 31433 63911 31467
rect 63911 31433 63920 31467
rect 63868 31424 63920 31433
rect 64144 31288 64196 31340
rect 77668 31331 77720 31340
rect 77668 31297 77677 31331
rect 77677 31297 77711 31331
rect 77711 31297 77720 31331
rect 77668 31288 77720 31297
rect 61844 31220 61896 31272
rect 61016 31152 61068 31204
rect 63040 31220 63092 31272
rect 62120 31084 62172 31136
rect 77852 31127 77904 31136
rect 77852 31093 77861 31127
rect 77861 31093 77895 31127
rect 77895 31093 77904 31127
rect 77852 31084 77904 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 62120 30787 62172 30796
rect 62120 30753 62129 30787
rect 62129 30753 62163 30787
rect 62163 30753 62172 30787
rect 62120 30744 62172 30753
rect 77668 30676 77720 30728
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 58440 30311 58492 30320
rect 58440 30277 58449 30311
rect 58449 30277 58483 30311
rect 58483 30277 58492 30311
rect 58440 30268 58492 30277
rect 58348 30132 58400 30184
rect 60464 30132 60516 30184
rect 61016 30064 61068 30116
rect 77852 30107 77904 30116
rect 77852 30073 77861 30107
rect 77861 30073 77895 30107
rect 77895 30073 77904 30107
rect 77852 30064 77904 30073
rect 58716 29996 58768 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 60464 29835 60516 29844
rect 60464 29801 60473 29835
rect 60473 29801 60507 29835
rect 60507 29801 60516 29835
rect 60464 29792 60516 29801
rect 58716 29699 58768 29708
rect 58716 29665 58725 29699
rect 58725 29665 58759 29699
rect 58759 29665 58768 29699
rect 58716 29656 58768 29665
rect 61016 29699 61068 29708
rect 61016 29665 61025 29699
rect 61025 29665 61059 29699
rect 61059 29665 61068 29699
rect 61016 29656 61068 29665
rect 60648 29520 60700 29572
rect 60740 29452 60792 29504
rect 78036 29495 78088 29504
rect 78036 29461 78045 29495
rect 78045 29461 78079 29495
rect 78079 29461 78088 29495
rect 78036 29452 78088 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 77852 28543 77904 28552
rect 77852 28509 77861 28543
rect 77861 28509 77895 28543
rect 77895 28509 77904 28543
rect 77852 28500 77904 28509
rect 78036 28407 78088 28416
rect 78036 28373 78045 28407
rect 78045 28373 78079 28407
rect 78079 28373 78088 28407
rect 78036 28364 78088 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 56324 28067 56376 28076
rect 56324 28033 56333 28067
rect 56333 28033 56367 28067
rect 56367 28033 56376 28067
rect 56324 28024 56376 28033
rect 77852 27820 77904 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 56324 27616 56376 27668
rect 52644 27480 52696 27532
rect 54392 27455 54444 27464
rect 54392 27421 54401 27455
rect 54401 27421 54435 27455
rect 54435 27421 54444 27455
rect 54392 27412 54444 27421
rect 56048 27455 56100 27464
rect 56048 27421 56057 27455
rect 56057 27421 56091 27455
rect 56091 27421 56100 27455
rect 56048 27412 56100 27421
rect 76196 27412 76248 27464
rect 54024 27319 54076 27328
rect 54024 27285 54033 27319
rect 54033 27285 54067 27319
rect 54067 27285 54076 27319
rect 54024 27276 54076 27285
rect 54576 27276 54628 27328
rect 56416 27276 56468 27328
rect 78036 27319 78088 27328
rect 78036 27285 78045 27319
rect 78045 27285 78079 27319
rect 78079 27285 78088 27319
rect 78036 27276 78088 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 54024 27004 54076 27056
rect 77668 26979 77720 26988
rect 77668 26945 77677 26979
rect 77677 26945 77711 26979
rect 77711 26945 77720 26979
rect 77668 26936 77720 26945
rect 76196 26732 76248 26784
rect 77852 26775 77904 26784
rect 77852 26741 77861 26775
rect 77861 26741 77895 26775
rect 77895 26741 77904 26775
rect 77852 26732 77904 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 50712 26392 50764 26444
rect 52644 26435 52696 26444
rect 52644 26401 52653 26435
rect 52653 26401 52687 26435
rect 52687 26401 52696 26435
rect 52644 26392 52696 26401
rect 52460 26367 52512 26376
rect 52460 26333 52469 26367
rect 52469 26333 52503 26367
rect 52503 26333 52512 26367
rect 52460 26324 52512 26333
rect 52920 26256 52972 26308
rect 77668 26256 77720 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 77668 25891 77720 25900
rect 77668 25857 77677 25891
rect 77677 25857 77711 25891
rect 77711 25857 77720 25891
rect 77668 25848 77720 25857
rect 77852 25687 77904 25696
rect 77852 25653 77861 25687
rect 77861 25653 77895 25687
rect 77895 25653 77904 25687
rect 77852 25644 77904 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 50712 25347 50764 25356
rect 50712 25313 50721 25347
rect 50721 25313 50755 25347
rect 50755 25313 50764 25347
rect 50712 25304 50764 25313
rect 50804 25236 50856 25288
rect 50712 25100 50764 25152
rect 77668 25100 77720 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 48872 24939 48924 24948
rect 48872 24905 48881 24939
rect 48881 24905 48915 24939
rect 48915 24905 48924 24939
rect 48872 24896 48924 24905
rect 49148 24760 49200 24812
rect 77668 24803 77720 24812
rect 77668 24769 77677 24803
rect 77677 24769 77711 24803
rect 77711 24769 77720 24803
rect 77668 24760 77720 24769
rect 49700 24692 49752 24744
rect 50620 24692 50672 24744
rect 49240 24556 49292 24608
rect 77852 24599 77904 24608
rect 77852 24565 77861 24599
rect 77861 24565 77895 24599
rect 77895 24565 77904 24599
rect 77852 24556 77904 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 49240 24191 49292 24200
rect 49240 24157 49249 24191
rect 49249 24157 49283 24191
rect 49283 24157 49292 24191
rect 49240 24148 49292 24157
rect 77668 24012 77720 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 49700 23851 49752 23860
rect 49700 23817 49709 23851
rect 49709 23817 49743 23851
rect 49743 23817 49752 23851
rect 49700 23808 49752 23817
rect 49608 23715 49660 23724
rect 49608 23681 49617 23715
rect 49617 23681 49651 23715
rect 49651 23681 49660 23715
rect 49608 23672 49660 23681
rect 47032 23604 47084 23656
rect 77852 23579 77904 23588
rect 77852 23545 77861 23579
rect 77861 23545 77895 23579
rect 77895 23545 77904 23579
rect 77852 23536 77904 23545
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 47032 23239 47084 23248
rect 47032 23205 47041 23239
rect 47041 23205 47075 23239
rect 47075 23205 47084 23239
rect 47032 23196 47084 23205
rect 46204 22992 46256 23044
rect 77484 22967 77536 22976
rect 77484 22933 77493 22967
rect 77493 22933 77527 22967
rect 77527 22933 77536 22967
rect 77484 22924 77536 22933
rect 78036 22967 78088 22976
rect 78036 22933 78045 22967
rect 78045 22933 78079 22967
rect 78079 22933 78088 22967
rect 78036 22924 78088 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 44824 22763 44876 22772
rect 44824 22729 44833 22763
rect 44833 22729 44867 22763
rect 44867 22729 44876 22763
rect 44824 22720 44876 22729
rect 46204 22763 46256 22772
rect 46204 22729 46213 22763
rect 46213 22729 46247 22763
rect 46247 22729 46256 22763
rect 46204 22720 46256 22729
rect 46572 22763 46624 22772
rect 46572 22729 46581 22763
rect 46581 22729 46615 22763
rect 46615 22729 46624 22763
rect 46572 22720 46624 22729
rect 45192 22652 45244 22704
rect 77484 22720 77536 22772
rect 45284 22584 45336 22636
rect 49976 22627 50028 22636
rect 49976 22593 49985 22627
rect 49985 22593 50019 22627
rect 50019 22593 50028 22627
rect 49976 22584 50028 22593
rect 46664 22559 46716 22568
rect 43168 22448 43220 22500
rect 46664 22525 46673 22559
rect 46673 22525 46707 22559
rect 46707 22525 46716 22559
rect 46664 22516 46716 22525
rect 45008 22380 45060 22432
rect 49608 22380 49660 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 45192 22219 45244 22228
rect 45192 22185 45201 22219
rect 45201 22185 45235 22219
rect 45235 22185 45244 22219
rect 45192 22176 45244 22185
rect 41696 22108 41748 22160
rect 43168 22108 43220 22160
rect 36544 21972 36596 22024
rect 42800 21972 42852 22024
rect 49608 22040 49660 22092
rect 45008 22015 45060 22024
rect 45008 21981 45017 22015
rect 45017 21981 45051 22015
rect 45051 21981 45060 22015
rect 45008 21972 45060 21981
rect 77852 22015 77904 22024
rect 77852 21981 77861 22015
rect 77861 21981 77895 22015
rect 77895 21981 77904 22015
rect 77852 21972 77904 21981
rect 43168 21836 43220 21888
rect 43904 21879 43956 21888
rect 43904 21845 43913 21879
rect 43913 21845 43947 21879
rect 43947 21845 43956 21879
rect 43904 21836 43956 21845
rect 78036 21879 78088 21888
rect 78036 21845 78045 21879
rect 78045 21845 78079 21879
rect 78079 21845 78088 21879
rect 78036 21836 78088 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 43904 21632 43956 21684
rect 77852 21632 77904 21684
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 41696 20995 41748 21004
rect 41696 20961 41705 20995
rect 41705 20961 41739 20995
rect 41739 20961 41748 20995
rect 41696 20952 41748 20961
rect 40224 20927 40276 20936
rect 40224 20893 40233 20927
rect 40233 20893 40267 20927
rect 40267 20893 40276 20927
rect 40224 20884 40276 20893
rect 41328 20884 41380 20936
rect 41604 20816 41656 20868
rect 39672 20748 39724 20800
rect 40132 20748 40184 20800
rect 41236 20748 41288 20800
rect 41512 20791 41564 20800
rect 41512 20757 41521 20791
rect 41521 20757 41555 20791
rect 41555 20757 41564 20791
rect 78036 20791 78088 20800
rect 41512 20748 41564 20757
rect 78036 20757 78045 20791
rect 78045 20757 78079 20791
rect 78079 20757 78088 20791
rect 78036 20748 78088 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 41604 20544 41656 20596
rect 39672 20451 39724 20460
rect 39672 20417 39681 20451
rect 39681 20417 39715 20451
rect 39715 20417 39724 20451
rect 39672 20408 39724 20417
rect 41236 20451 41288 20460
rect 41236 20417 41245 20451
rect 41245 20417 41279 20451
rect 41279 20417 41288 20451
rect 41236 20408 41288 20417
rect 49976 20408 50028 20460
rect 50988 20383 51040 20392
rect 50988 20349 50997 20383
rect 50997 20349 51031 20383
rect 51031 20349 51040 20383
rect 50988 20340 51040 20349
rect 77116 20340 77168 20392
rect 77852 20247 77904 20256
rect 77852 20213 77861 20247
rect 77861 20213 77895 20247
rect 77895 20213 77904 20247
rect 77852 20204 77904 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 77300 19320 77352 19372
rect 77300 19159 77352 19168
rect 77300 19125 77309 19159
rect 77309 19125 77343 19159
rect 77343 19125 77352 19159
rect 77300 19116 77352 19125
rect 77852 19159 77904 19168
rect 77852 19125 77861 19159
rect 77861 19125 77895 19159
rect 77895 19125 77904 19159
rect 77852 19116 77904 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 37280 18708 37332 18760
rect 77300 18572 77352 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 37280 18411 37332 18420
rect 37280 18377 37289 18411
rect 37289 18377 37323 18411
rect 37323 18377 37332 18411
rect 37280 18368 37332 18377
rect 37648 18411 37700 18420
rect 37648 18377 37657 18411
rect 37657 18377 37691 18411
rect 37691 18377 37700 18411
rect 37648 18368 37700 18377
rect 36268 18232 36320 18284
rect 37556 18164 37608 18216
rect 36728 18096 36780 18148
rect 77852 18071 77904 18080
rect 77852 18037 77861 18071
rect 77861 18037 77895 18071
rect 77895 18037 77904 18071
rect 77852 18028 77904 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 36268 17867 36320 17876
rect 36268 17833 36277 17867
rect 36277 17833 36311 17867
rect 36311 17833 36320 17867
rect 36268 17824 36320 17833
rect 33692 17688 33744 17740
rect 35440 17552 35492 17604
rect 77852 17663 77904 17672
rect 77852 17629 77861 17663
rect 77861 17629 77895 17663
rect 77895 17629 77904 17663
rect 77852 17620 77904 17629
rect 36728 17552 36780 17604
rect 35532 17484 35584 17536
rect 78036 17527 78088 17536
rect 78036 17493 78045 17527
rect 78045 17493 78079 17527
rect 78079 17493 78088 17527
rect 78036 17484 78088 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 33324 17280 33376 17332
rect 31668 17212 31720 17264
rect 33692 17212 33744 17264
rect 36544 17255 36596 17264
rect 36544 17221 36553 17255
rect 36553 17221 36587 17255
rect 36587 17221 36596 17255
rect 36544 17212 36596 17221
rect 36728 17255 36780 17264
rect 36728 17221 36737 17255
rect 36737 17221 36771 17255
rect 36771 17221 36780 17255
rect 36728 17212 36780 17221
rect 33508 17119 33560 17128
rect 33508 17085 33517 17119
rect 33517 17085 33551 17119
rect 33551 17085 33560 17119
rect 33508 17076 33560 17085
rect 77852 16940 77904 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 31576 16643 31628 16652
rect 31576 16609 31585 16643
rect 31585 16609 31619 16643
rect 31619 16609 31628 16643
rect 31576 16600 31628 16609
rect 31668 16643 31720 16652
rect 31668 16609 31677 16643
rect 31677 16609 31711 16643
rect 31711 16609 31720 16643
rect 31668 16600 31720 16609
rect 32404 16532 32456 16584
rect 77852 16575 77904 16584
rect 77852 16541 77861 16575
rect 77861 16541 77895 16575
rect 77895 16541 77904 16575
rect 77852 16532 77904 16541
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 78036 16439 78088 16448
rect 78036 16405 78045 16439
rect 78045 16405 78079 16439
rect 78079 16405 78088 16439
rect 78036 16396 78088 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 29920 16235 29972 16244
rect 29920 16201 29929 16235
rect 29929 16201 29963 16235
rect 29963 16201 29972 16235
rect 29920 16192 29972 16201
rect 31116 16124 31168 16176
rect 29552 15988 29604 16040
rect 31668 15988 31720 16040
rect 30288 15852 30340 15904
rect 77852 15852 77904 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 12440 15648 12492 15700
rect 30288 15487 30340 15496
rect 30288 15453 30297 15487
rect 30297 15453 30331 15487
rect 30331 15453 30340 15487
rect 30288 15444 30340 15453
rect 14280 15419 14332 15428
rect 14280 15385 14289 15419
rect 14289 15385 14323 15419
rect 14323 15385 14332 15419
rect 14280 15376 14332 15385
rect 78036 15351 78088 15360
rect 78036 15317 78045 15351
rect 78045 15317 78079 15351
rect 78079 15317 78088 15351
rect 78036 15308 78088 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 16764 15104 16816 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 14648 14968 14700 15020
rect 16304 14968 16356 15020
rect 17776 14968 17828 15020
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 14372 14900 14424 14952
rect 1400 14764 1452 14816
rect 15384 14764 15436 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 14280 14560 14332 14612
rect 16304 14603 16356 14612
rect 16304 14569 16313 14603
rect 16313 14569 16347 14603
rect 16347 14569 16356 14603
rect 16304 14560 16356 14569
rect 14004 14492 14056 14544
rect 16212 14535 16264 14544
rect 16212 14501 16221 14535
rect 16221 14501 16255 14535
rect 16255 14501 16264 14535
rect 16212 14492 16264 14501
rect 17684 14492 17736 14544
rect 14188 14331 14240 14340
rect 14188 14297 14197 14331
rect 14197 14297 14231 14331
rect 14231 14297 14240 14331
rect 14188 14288 14240 14297
rect 17776 14220 17828 14272
rect 27252 14288 27304 14340
rect 36544 14288 36596 14340
rect 27160 14263 27212 14272
rect 27160 14229 27169 14263
rect 27169 14229 27203 14263
rect 27203 14229 27212 14263
rect 27160 14220 27212 14229
rect 78036 14263 78088 14272
rect 78036 14229 78045 14263
rect 78045 14229 78079 14263
rect 78079 14229 78088 14263
rect 78036 14220 78088 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 27252 14016 27304 14068
rect 27528 14059 27580 14068
rect 27528 14025 27537 14059
rect 27537 14025 27571 14059
rect 27571 14025 27580 14059
rect 27528 14016 27580 14025
rect 14188 13991 14240 14000
rect 14188 13957 14197 13991
rect 14197 13957 14231 13991
rect 14231 13957 14240 13991
rect 14188 13948 14240 13957
rect 26976 13948 27028 14000
rect 27344 13812 27396 13864
rect 14464 13787 14516 13796
rect 14464 13753 14473 13787
rect 14473 13753 14507 13787
rect 14507 13753 14516 13787
rect 14464 13744 14516 13753
rect 27160 13744 27212 13796
rect 77852 13719 77904 13728
rect 77852 13685 77861 13719
rect 77861 13685 77895 13719
rect 77895 13685 77904 13719
rect 77852 13676 77904 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 26976 13515 27028 13524
rect 26976 13481 26985 13515
rect 26985 13481 27019 13515
rect 27019 13481 27028 13515
rect 26976 13472 27028 13481
rect 25964 13379 26016 13388
rect 25964 13345 25973 13379
rect 25973 13345 26007 13379
rect 26007 13345 26016 13379
rect 25964 13336 26016 13345
rect 27160 13336 27212 13388
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 25688 13132 25740 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 24768 12588 24820 12640
rect 77852 12631 77904 12640
rect 77852 12597 77861 12631
rect 77861 12597 77895 12631
rect 77895 12597 77904 12631
rect 77852 12588 77904 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 24768 12427 24820 12436
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 23664 12291 23716 12300
rect 23664 12257 23673 12291
rect 23673 12257 23707 12291
rect 23707 12257 23716 12291
rect 23664 12248 23716 12257
rect 25964 12248 26016 12300
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 23480 12180 23532 12189
rect 24400 12044 24452 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 22192 11883 22244 11892
rect 22192 11849 22201 11883
rect 22201 11849 22235 11883
rect 22235 11849 22244 11883
rect 22192 11840 22244 11849
rect 20076 11636 20128 11688
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 23664 11636 23716 11688
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 77852 11611 77904 11620
rect 77852 11577 77861 11611
rect 77861 11577 77895 11611
rect 77895 11577 77904 11611
rect 77852 11568 77904 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 78036 11271 78088 11280
rect 78036 11237 78045 11271
rect 78045 11237 78079 11271
rect 78079 11237 78088 11271
rect 78036 11228 78088 11237
rect 19984 11092 20036 11144
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 77944 10115 77996 10124
rect 77944 10081 77953 10115
rect 77953 10081 77987 10115
rect 77987 10081 77996 10115
rect 77944 10072 77996 10081
rect 77668 10047 77720 10056
rect 77668 10013 77677 10047
rect 77677 10013 77711 10047
rect 77711 10013 77720 10047
rect 77668 10004 77720 10013
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 2872 9052 2924 9104
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 77668 8959 77720 8968
rect 77668 8925 77677 8959
rect 77677 8925 77711 8959
rect 77711 8925 77720 8959
rect 77668 8916 77720 8925
rect 8392 8848 8444 8900
rect 77576 8848 77628 8900
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4804 8576 4856 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 9036 8440 9088 8492
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 6736 8304 6788 8356
rect 10048 8304 10100 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 8944 8032 8996 8084
rect 10508 8032 10560 8084
rect 9128 7964 9180 8016
rect 9312 8007 9364 8016
rect 9312 7973 9321 8007
rect 9321 7973 9355 8007
rect 9355 7973 9364 8007
rect 9312 7964 9364 7973
rect 10324 7896 10376 7948
rect 77668 7871 77720 7880
rect 77668 7837 77677 7871
rect 77677 7837 77711 7871
rect 77711 7837 77720 7871
rect 77668 7828 77720 7837
rect 8760 7760 8812 7812
rect 78036 7760 78088 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 9036 7488 9088 7540
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 9956 7352 10008 7404
rect 77208 7352 77260 7404
rect 77852 7284 77904 7336
rect 9404 7216 9456 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 77484 6307 77536 6316
rect 77484 6273 77493 6307
rect 77493 6273 77527 6307
rect 77527 6273 77536 6307
rect 77484 6264 77536 6273
rect 77392 6196 77444 6248
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 77484 5219 77536 5228
rect 77484 5185 77493 5219
rect 77493 5185 77527 5219
rect 77527 5185 77536 5219
rect 77484 5176 77536 5185
rect 77484 4972 77536 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 77668 4607 77720 4616
rect 77668 4573 77677 4607
rect 77677 4573 77711 4607
rect 77711 4573 77720 4607
rect 77668 4564 77720 4573
rect 77300 4496 77352 4548
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 79048 4156 79100 4208
rect 9128 4088 9180 4140
rect 9588 4088 9640 4140
rect 77300 4088 77352 4140
rect 78128 4088 78180 4140
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 9588 3723 9640 3732
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 14004 3612 14056 3664
rect 21364 3612 21416 3664
rect 9680 3544 9732 3596
rect 77760 3544 77812 3596
rect 9956 3519 10008 3528
rect 8116 3340 8168 3392
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 14372 3476 14424 3528
rect 16672 3476 16724 3528
rect 50988 3476 51040 3528
rect 77668 3519 77720 3528
rect 77668 3485 77677 3519
rect 77677 3485 77711 3519
rect 77711 3485 77720 3519
rect 77668 3476 77720 3485
rect 21364 3408 21416 3460
rect 77392 3408 77444 3460
rect 77944 3451 77996 3460
rect 77944 3417 77953 3451
rect 77953 3417 77987 3451
rect 77987 3417 77996 3451
rect 77944 3408 77996 3417
rect 9864 3340 9916 3392
rect 13820 3340 13872 3392
rect 15108 3340 15160 3392
rect 16580 3340 16632 3392
rect 76288 3340 76340 3392
rect 78036 3340 78088 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16672 3179 16724 3188
rect 16212 3136 16264 3145
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 14280 3000 14332 3052
rect 14648 3000 14700 3052
rect 15108 3000 15160 3052
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 76288 3136 76340 3188
rect 76932 3179 76984 3188
rect 76932 3145 76941 3179
rect 76941 3145 76975 3179
rect 76975 3145 76984 3179
rect 76932 3136 76984 3145
rect 15384 3000 15436 3009
rect 7564 2864 7616 2916
rect 15108 2864 15160 2916
rect 77944 3068 77996 3120
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 41512 3000 41564 3052
rect 77116 3000 77168 3052
rect 77760 3043 77812 3052
rect 40960 2932 41012 2984
rect 77024 2932 77076 2984
rect 77760 3009 77769 3043
rect 77769 3009 77803 3043
rect 77803 3009 77812 3043
rect 77760 3000 77812 3009
rect 77576 2864 77628 2916
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 8392 2796 8444 2848
rect 14096 2796 14148 2848
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 20076 2635 20128 2644
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 22284 2592 22336 2644
rect 24400 2635 24452 2644
rect 24400 2601 24409 2635
rect 24409 2601 24443 2635
rect 24443 2601 24452 2635
rect 24400 2592 24452 2601
rect 25688 2592 25740 2644
rect 27344 2592 27396 2644
rect 29552 2635 29604 2644
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 29552 2592 29604 2601
rect 31576 2592 31628 2644
rect 46664 2592 46716 2644
rect 49148 2592 49200 2644
rect 50712 2635 50764 2644
rect 50712 2601 50721 2635
rect 50721 2601 50755 2635
rect 50755 2601 50764 2635
rect 50712 2592 50764 2601
rect 52920 2635 52972 2644
rect 52920 2601 52929 2635
rect 52929 2601 52963 2635
rect 52963 2601 52972 2635
rect 52920 2592 52972 2601
rect 54576 2635 54628 2644
rect 54576 2601 54585 2635
rect 54585 2601 54619 2635
rect 54619 2601 54628 2635
rect 54576 2592 54628 2601
rect 56416 2635 56468 2644
rect 56416 2601 56425 2635
rect 56425 2601 56459 2635
rect 56459 2601 56468 2635
rect 56416 2592 56468 2601
rect 58348 2635 58400 2644
rect 58348 2601 58357 2635
rect 58357 2601 58391 2635
rect 58391 2601 58400 2635
rect 58348 2592 58400 2601
rect 61844 2592 61896 2644
rect 64144 2592 64196 2644
rect 66076 2592 66128 2644
rect 68376 2635 68428 2644
rect 68376 2601 68385 2635
rect 68385 2601 68419 2635
rect 68419 2601 68428 2635
rect 68376 2592 68428 2601
rect 69848 2592 69900 2644
rect 71412 2592 71464 2644
rect 73620 2635 73672 2644
rect 73620 2601 73629 2635
rect 73629 2601 73663 2635
rect 73663 2601 73672 2635
rect 73620 2592 73672 2601
rect 75184 2592 75236 2644
rect 7564 2388 7616 2440
rect 8392 2456 8444 2508
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10324 2388 10376 2440
rect 13820 2456 13872 2508
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 8208 2320 8260 2372
rect 940 2252 992 2304
rect 2780 2252 2832 2304
rect 4712 2252 4764 2304
rect 6644 2252 6696 2304
rect 8484 2252 8536 2304
rect 10416 2252 10468 2304
rect 14096 2388 14148 2440
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 77852 2524 77904 2576
rect 15384 2456 15436 2508
rect 14464 2388 14516 2397
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 16580 2388 16632 2440
rect 18328 2388 18380 2440
rect 19984 2388 20036 2440
rect 21824 2388 21876 2440
rect 23756 2388 23808 2440
rect 25688 2388 25740 2440
rect 27620 2388 27672 2440
rect 29460 2388 29512 2440
rect 31392 2388 31444 2440
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 33508 2388 33560 2440
rect 35164 2388 35216 2440
rect 35532 2431 35584 2440
rect 35532 2397 35541 2431
rect 35541 2397 35575 2431
rect 35575 2397 35584 2431
rect 35532 2388 35584 2397
rect 37096 2388 37148 2440
rect 37556 2431 37608 2440
rect 37556 2397 37565 2431
rect 37565 2397 37599 2431
rect 37599 2397 37608 2431
rect 37556 2388 37608 2397
rect 39028 2388 39080 2440
rect 40132 2431 40184 2440
rect 40132 2397 40141 2431
rect 40141 2397 40175 2431
rect 40175 2397 40184 2431
rect 40132 2388 40184 2397
rect 42800 2388 42852 2440
rect 43168 2431 43220 2440
rect 43168 2397 43177 2431
rect 43177 2397 43211 2431
rect 43211 2397 43220 2431
rect 43168 2388 43220 2397
rect 44732 2388 44784 2440
rect 45284 2431 45336 2440
rect 45284 2397 45293 2431
rect 45293 2397 45327 2431
rect 45327 2397 45336 2431
rect 45284 2388 45336 2397
rect 46664 2388 46716 2440
rect 60740 2431 60792 2440
rect 60740 2397 60749 2431
rect 60749 2397 60783 2431
rect 60783 2397 60792 2431
rect 60740 2388 60792 2397
rect 73344 2388 73396 2440
rect 75184 2388 75236 2440
rect 76564 2431 76616 2440
rect 76564 2397 76573 2431
rect 76573 2397 76607 2431
rect 76607 2397 76616 2431
rect 76564 2388 76616 2397
rect 77208 2388 77260 2440
rect 14280 2320 14332 2372
rect 12348 2252 12400 2304
rect 48504 2320 48556 2372
rect 50620 2363 50672 2372
rect 50620 2329 50629 2363
rect 50629 2329 50663 2363
rect 50663 2329 50672 2363
rect 50620 2320 50672 2329
rect 52368 2320 52420 2372
rect 54300 2320 54352 2372
rect 56140 2320 56192 2372
rect 58072 2320 58124 2372
rect 60004 2320 60056 2372
rect 61844 2320 61896 2372
rect 63776 2320 63828 2372
rect 65708 2320 65760 2372
rect 67640 2320 67692 2372
rect 69480 2320 69532 2372
rect 71412 2320 71464 2372
rect 77760 2363 77812 2372
rect 77760 2329 77769 2363
rect 77769 2329 77803 2363
rect 77803 2329 77812 2363
rect 77760 2320 77812 2329
rect 16120 2252 16172 2304
rect 18052 2252 18104 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 9956 1980 10008 2032
rect 77484 1980 77536 2032
rect 9128 1912 9180 1964
rect 77760 1912 77812 1964
<< metal2 >>
rect 938 39200 994 40000
rect 2778 39200 2834 40000
rect 4710 39200 4766 40000
rect 6642 39200 6698 40000
rect 8482 39200 8538 40000
rect 10414 39200 10470 40000
rect 12346 39200 12402 40000
rect 14278 39200 14334 40000
rect 16118 39200 16174 40000
rect 16224 39222 16528 39250
rect 952 37126 980 39200
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 940 37120 992 37126
rect 940 37062 992 37068
rect 1412 14822 1440 37198
rect 2792 37126 2820 39200
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 2872 37256 2924 37262
rect 2872 37198 2924 37204
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 2884 9110 2912 37198
rect 4724 37126 4752 39200
rect 4804 37256 4856 37262
rect 4804 37198 4856 37204
rect 4712 37120 4764 37126
rect 4712 37062 4764 37068
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 4816 8634 4844 37198
rect 6656 37126 6684 39200
rect 6736 37256 6788 37262
rect 6736 37198 6788 37204
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 6644 37120 6696 37126
rect 6644 37062 6696 37068
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 6748 8362 6776 37198
rect 8312 9178 8340 37198
rect 8496 37126 8524 39200
rect 10428 37126 10456 39200
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 8484 37120 8536 37126
rect 8484 37062 8536 37068
rect 10416 37120 10468 37126
rect 10416 37062 10468 37068
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 8404 8090 8432 8842
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8772 7818 8800 8366
rect 8956 8090 8984 8910
rect 10612 8634 10640 37198
rect 12360 37126 12388 39200
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 12452 15706 12480 37198
rect 14292 37126 14320 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 16500 37210 16528 39222
rect 18050 39200 18106 40000
rect 19982 39200 20038 40000
rect 21822 39200 21878 40000
rect 23754 39200 23810 40000
rect 25686 39200 25742 40000
rect 27618 39200 27674 40000
rect 29458 39200 29514 40000
rect 31390 39200 31446 40000
rect 33322 39200 33378 40000
rect 35162 39200 35218 40000
rect 37094 39200 37150 40000
rect 39026 39200 39082 40000
rect 40958 39200 41014 40000
rect 42798 39200 42854 40000
rect 44730 39200 44786 40000
rect 46662 39200 46718 40000
rect 48502 39200 48558 40000
rect 50434 39200 50490 40000
rect 52366 39200 52422 40000
rect 54298 39200 54354 40000
rect 56138 39200 56194 40000
rect 58070 39200 58126 40000
rect 60002 39200 60058 40000
rect 61842 39200 61898 40000
rect 63774 39200 63830 40000
rect 65706 39200 65762 40000
rect 65812 39222 66024 39250
rect 16764 37256 16816 37262
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8772 7478 8800 7754
rect 9048 7546 9076 8434
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 9140 4146 9168 7958
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9324 4026 9352 7958
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9140 3998 9352 4026
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 7576 2446 7604 2858
rect 8128 2446 8156 3334
rect 9140 3058 9168 3998
rect 9416 3618 9444 7210
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3738 9628 4082
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9416 3602 9720 3618
rect 9416 3596 9732 3602
rect 9416 3590 9680 3596
rect 9600 3058 9628 3590
rect 9680 3538 9732 3544
rect 9968 3534 9996 7346
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8220 2378 8248 2790
rect 8404 2514 8432 2790
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 952 800 980 2246
rect 2792 800 2820 2246
rect 4724 800 4752 2246
rect 6656 800 6684 2246
rect 8496 800 8524 2246
rect 9140 1970 9168 2994
rect 9876 2990 9904 3334
rect 10060 3058 10088 8298
rect 10520 8090 10548 8434
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9876 2446 9904 2926
rect 10336 2446 10364 7890
rect 14016 3670 14044 14486
rect 14200 14346 14228 14894
rect 14292 14618 14320 15370
rect 14384 14958 14412 37198
rect 16500 37182 16620 37210
rect 16764 37198 16816 37204
rect 16592 37126 16620 37182
rect 16580 37120 16632 37126
rect 16580 37062 16632 37068
rect 16776 15162 16804 37198
rect 18064 37126 18092 39200
rect 19996 37262 20024 39200
rect 20352 37324 20404 37330
rect 20352 37266 20404 37272
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18432 15162 18460 37198
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14200 14006 14228 14282
rect 14660 14074 14688 14962
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13832 2514 13860 3334
rect 14016 3194 14044 3606
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3194 14412 3470
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14108 2446 14136 2790
rect 14292 2650 14320 2994
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14476 2446 14504 13738
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15120 3058 15148 3334
rect 15396 3058 15424 14758
rect 16316 14618 16344 14962
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 16224 3194 16252 14486
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 14660 2514 14688 2994
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15120 2446 15148 2858
rect 15396 2514 15424 2994
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 16592 2446 16620 3334
rect 16684 3194 16712 3470
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17696 3058 17724 14486
rect 17788 14278 17816 14962
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20364 11898 20392 37266
rect 21836 37262 21864 39200
rect 22192 37324 22244 37330
rect 22192 37266 22244 37272
rect 23480 37324 23532 37330
rect 23480 37266 23532 37272
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 22204 11898 22232 37266
rect 23492 12238 23520 37266
rect 23768 37262 23796 39200
rect 25700 37262 25728 39200
rect 25780 37324 25832 37330
rect 25780 37266 25832 37272
rect 27528 37324 27580 37330
rect 27528 37266 27580 37272
rect 23756 37256 23808 37262
rect 23756 37198 23808 37204
rect 25688 37256 25740 37262
rect 25688 37198 25740 37204
rect 25792 13326 25820 37266
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 26976 14000 27028 14006
rect 26976 13942 27028 13948
rect 26988 13530 27016 13942
rect 27172 13802 27200 14214
rect 27264 14074 27292 14282
rect 27540 14074 27568 37266
rect 27632 37262 27660 39200
rect 29472 37330 29500 39200
rect 31404 37330 31432 39200
rect 29460 37324 29512 37330
rect 29460 37266 29512 37272
rect 31392 37324 31444 37330
rect 31392 37266 31444 37272
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 29920 37256 29972 37262
rect 29920 37198 29972 37204
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 29932 16250 29960 37198
rect 31668 17264 31720 17270
rect 31668 17206 31720 17212
rect 31680 16658 31708 17206
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31668 16652 31720 16658
rect 31668 16594 31720 16600
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 31128 16182 31156 16390
rect 31116 16176 31168 16182
rect 31116 16118 31168 16124
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27172 13394 27200 13738
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24780 12442 24808 12582
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 23676 11694 23704 12242
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11150 20024 11494
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2446 18368 2790
rect 20088 2650 20116 11630
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21376 3466 21404 3606
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 22296 2650 22324 11630
rect 24412 2650 24440 12038
rect 25700 2650 25728 13126
rect 25976 12306 26004 13330
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 27356 2650 27384 13806
rect 29564 2650 29592 15982
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30300 15502 30328 15846
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 31588 2650 31616 16594
rect 31680 16046 31708 16594
rect 32416 16590 32444 37198
rect 33336 36786 33364 39200
rect 35176 38298 35204 39200
rect 35176 38270 35388 38298
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35360 37330 35388 38270
rect 37108 37330 37136 39200
rect 39040 37330 39068 39200
rect 35348 37324 35400 37330
rect 35348 37266 35400 37272
rect 37096 37324 37148 37330
rect 37096 37266 37148 37272
rect 39028 37324 39080 37330
rect 39028 37266 39080 37272
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 37648 37256 37700 37262
rect 37648 37198 37700 37204
rect 40224 37256 40276 37262
rect 40224 37198 40276 37204
rect 33324 36780 33376 36786
rect 33324 36722 33376 36728
rect 33324 36644 33376 36650
rect 33324 36586 33376 36592
rect 33336 17338 33364 36586
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 33692 17740 33744 17746
rect 33692 17682 33744 17688
rect 33324 17332 33376 17338
rect 33324 17274 33376 17280
rect 33704 17270 33732 17682
rect 35452 17610 35480 37198
rect 36544 22024 36596 22030
rect 36544 21966 36596 21972
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36280 17882 36308 18226
rect 36268 17876 36320 17882
rect 36268 17818 36320 17824
rect 35440 17604 35492 17610
rect 35440 17546 35492 17552
rect 35532 17536 35584 17542
rect 35532 17478 35584 17484
rect 33692 17264 33744 17270
rect 33692 17206 33744 17212
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 31668 16040 31720 16046
rect 31668 15982 31720 15988
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 31576 2644 31628 2650
rect 31576 2586 31628 2592
rect 33520 2446 33548 17070
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35544 2446 35572 17478
rect 36556 17270 36584 21966
rect 37280 18760 37332 18766
rect 37280 18702 37332 18708
rect 37292 18426 37320 18702
rect 37660 18426 37688 37198
rect 40236 20942 40264 37198
rect 40972 36786 41000 39200
rect 42812 37330 42840 39200
rect 44744 37330 44772 39200
rect 42800 37324 42852 37330
rect 42800 37266 42852 37272
rect 44732 37324 44784 37330
rect 44732 37266 44784 37272
rect 46676 37262 46704 39200
rect 48516 37262 48544 39200
rect 50448 37262 50476 39200
rect 44824 37256 44876 37262
rect 44824 37198 44876 37204
rect 46664 37256 46716 37262
rect 46664 37198 46716 37204
rect 48504 37256 48556 37262
rect 48504 37198 48556 37204
rect 50436 37256 50488 37262
rect 50436 37198 50488 37204
rect 52380 37210 52408 39200
rect 54312 37262 54340 39200
rect 56152 37262 56180 39200
rect 58084 37262 58112 39200
rect 60016 37262 60044 39200
rect 61856 37262 61884 39200
rect 63788 37262 63816 39200
rect 65720 39114 65748 39200
rect 65812 39114 65840 39222
rect 65720 39086 65840 39114
rect 65654 37564 65962 37584
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37488 65962 37508
rect 65996 37262 66024 39222
rect 67638 39200 67694 40000
rect 69478 39200 69534 40000
rect 71410 39200 71466 40000
rect 73342 39200 73398 40000
rect 75182 39200 75238 40000
rect 76746 39536 76802 39545
rect 76746 39471 76802 39480
rect 67652 37262 67680 39200
rect 69492 37262 69520 39200
rect 71424 37262 71452 39200
rect 73356 37262 73384 39200
rect 75196 37262 75224 39200
rect 52460 37256 52512 37262
rect 52380 37204 52460 37210
rect 52380 37198 52512 37204
rect 54300 37256 54352 37262
rect 54300 37198 54352 37204
rect 56140 37256 56192 37262
rect 56140 37198 56192 37204
rect 58072 37256 58124 37262
rect 58072 37198 58124 37204
rect 60004 37256 60056 37262
rect 60004 37198 60056 37204
rect 61844 37256 61896 37262
rect 61844 37198 61896 37204
rect 63776 37256 63828 37262
rect 63776 37198 63828 37204
rect 65984 37256 66036 37262
rect 65984 37198 66036 37204
rect 67640 37256 67692 37262
rect 67640 37198 67692 37204
rect 69480 37256 69532 37262
rect 69480 37198 69532 37204
rect 71412 37256 71464 37262
rect 71412 37198 71464 37204
rect 73344 37256 73396 37262
rect 73344 37198 73396 37204
rect 75184 37256 75236 37262
rect 75184 37198 75236 37204
rect 42800 37188 42852 37194
rect 42800 37130 42852 37136
rect 40960 36780 41012 36786
rect 40960 36722 41012 36728
rect 41328 36712 41380 36718
rect 41328 36654 41380 36660
rect 41340 20942 41368 36654
rect 41696 22160 41748 22166
rect 41696 22102 41748 22108
rect 41708 21010 41736 22102
rect 42812 22030 42840 37130
rect 44836 22778 44864 37198
rect 52380 37182 52500 37198
rect 74724 37188 74776 37194
rect 74724 37130 74776 37136
rect 46572 37120 46624 37126
rect 46572 37062 46624 37068
rect 48872 37120 48924 37126
rect 48872 37062 48924 37068
rect 50804 37120 50856 37126
rect 50804 37062 50856 37068
rect 52460 37120 52512 37126
rect 52460 37062 52512 37068
rect 54392 37120 54444 37126
rect 54392 37062 54444 37068
rect 56048 37120 56100 37126
rect 56048 37062 56100 37068
rect 58440 37120 58492 37126
rect 58440 37062 58492 37068
rect 60648 37120 60700 37126
rect 60648 37062 60700 37068
rect 61936 37120 61988 37126
rect 61936 37062 61988 37068
rect 63868 37120 63920 37126
rect 63868 37062 63920 37068
rect 66168 37120 66220 37126
rect 66168 37062 66220 37068
rect 68192 37120 68244 37126
rect 68192 37062 68244 37068
rect 69572 37120 69624 37126
rect 69572 37062 69624 37068
rect 71504 37120 71556 37126
rect 71504 37062 71556 37068
rect 73712 37120 73764 37126
rect 73712 37062 73764 37068
rect 46204 23044 46256 23050
rect 46204 22986 46256 22992
rect 46216 22778 46244 22986
rect 46584 22778 46612 37062
rect 48884 24954 48912 37062
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 49976 31816 50028 31822
rect 49976 31758 50028 31764
rect 48872 24948 48924 24954
rect 48872 24890 48924 24896
rect 49148 24812 49200 24818
rect 49148 24754 49200 24760
rect 47032 23656 47084 23662
rect 47032 23598 47084 23604
rect 47044 23254 47072 23598
rect 47032 23248 47084 23254
rect 47032 23190 47084 23196
rect 44824 22772 44876 22778
rect 44824 22714 44876 22720
rect 46204 22772 46256 22778
rect 46204 22714 46256 22720
rect 46572 22772 46624 22778
rect 46572 22714 46624 22720
rect 45192 22704 45244 22710
rect 45192 22646 45244 22652
rect 43168 22500 43220 22506
rect 43168 22442 43220 22448
rect 43180 22166 43208 22442
rect 45008 22432 45060 22438
rect 45008 22374 45060 22380
rect 43168 22160 43220 22166
rect 43168 22102 43220 22108
rect 45020 22030 45048 22374
rect 45204 22234 45232 22646
rect 45284 22636 45336 22642
rect 45284 22578 45336 22584
rect 45192 22228 45244 22234
rect 45192 22170 45244 22176
rect 42800 22024 42852 22030
rect 42800 21966 42852 21972
rect 45008 22024 45060 22030
rect 45008 21966 45060 21972
rect 43168 21888 43220 21894
rect 43168 21830 43220 21836
rect 43904 21888 43956 21894
rect 43904 21830 43956 21836
rect 41696 21004 41748 21010
rect 41696 20946 41748 20952
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 41328 20936 41380 20942
rect 41328 20878 41380 20884
rect 41604 20868 41656 20874
rect 41604 20810 41656 20816
rect 39672 20800 39724 20806
rect 39672 20742 39724 20748
rect 40132 20800 40184 20806
rect 40132 20742 40184 20748
rect 41236 20800 41288 20806
rect 41236 20742 41288 20748
rect 41512 20800 41564 20806
rect 41512 20742 41564 20748
rect 39684 20466 39712 20742
rect 39672 20460 39724 20466
rect 39672 20402 39724 20408
rect 37280 18420 37332 18426
rect 37280 18362 37332 18368
rect 37648 18420 37700 18426
rect 37648 18362 37700 18368
rect 37556 18216 37608 18222
rect 37556 18158 37608 18164
rect 36728 18148 36780 18154
rect 36728 18090 36780 18096
rect 36740 17610 36768 18090
rect 36728 17604 36780 17610
rect 36728 17546 36780 17552
rect 36740 17270 36768 17546
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36728 17264 36780 17270
rect 36728 17206 36780 17212
rect 36556 14346 36584 17206
rect 36544 14340 36596 14346
rect 36544 14282 36596 14288
rect 37568 2446 37596 18158
rect 40144 2446 40172 20742
rect 41248 20466 41276 20742
rect 41236 20460 41288 20466
rect 41236 20402 41288 20408
rect 41524 3058 41552 20742
rect 41616 20602 41644 20810
rect 41604 20596 41656 20602
rect 41604 20538 41656 20544
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 40960 2984 41012 2990
rect 40960 2926 41012 2932
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 39028 2440 39080 2446
rect 39028 2382 39080 2388
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 9968 2038 9996 2382
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 9956 2032 10008 2038
rect 9956 1974 10008 1980
rect 9128 1964 9180 1970
rect 9128 1906 9180 1912
rect 10428 800 10456 2246
rect 12360 800 12388 2246
rect 14292 800 14320 2314
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 16132 800 16160 2246
rect 18064 800 18092 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2382
rect 21836 800 21864 2382
rect 23768 800 23796 2382
rect 25700 800 25728 2382
rect 27632 800 27660 2382
rect 29472 800 29500 2382
rect 31404 800 31432 2382
rect 33336 800 33364 2382
rect 35176 800 35204 2382
rect 37108 800 37136 2382
rect 39040 800 39068 2382
rect 40972 800 41000 2926
rect 43180 2446 43208 21830
rect 43916 21690 43944 21830
rect 43904 21684 43956 21690
rect 43904 21626 43956 21632
rect 45296 2446 45324 22578
rect 46664 22568 46716 22574
rect 46664 22510 46716 22516
rect 46676 2650 46704 22510
rect 49160 2650 49188 24754
rect 49700 24744 49752 24750
rect 49700 24686 49752 24692
rect 49240 24608 49292 24614
rect 49240 24550 49292 24556
rect 49252 24206 49280 24550
rect 49240 24200 49292 24206
rect 49240 24142 49292 24148
rect 49712 23866 49740 24686
rect 49700 23860 49752 23866
rect 49700 23802 49752 23808
rect 49608 23724 49660 23730
rect 49608 23666 49660 23672
rect 49620 22438 49648 23666
rect 49988 22642 50016 31758
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50712 26444 50764 26450
rect 50712 26386 50764 26392
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50724 25362 50752 26386
rect 50712 25356 50764 25362
rect 50712 25298 50764 25304
rect 50724 25242 50752 25298
rect 50816 25294 50844 37062
rect 52472 26382 52500 37062
rect 52644 27532 52696 27538
rect 52644 27474 52696 27480
rect 52656 26450 52684 27474
rect 54404 27470 54432 37062
rect 56060 27470 56088 37062
rect 58452 30326 58480 37062
rect 58440 30320 58492 30326
rect 58440 30262 58492 30268
rect 58348 30184 58400 30190
rect 58348 30126 58400 30132
rect 60464 30184 60516 30190
rect 60464 30126 60516 30132
rect 56324 28076 56376 28082
rect 56324 28018 56376 28024
rect 56336 27674 56364 28018
rect 56324 27668 56376 27674
rect 56324 27610 56376 27616
rect 54392 27464 54444 27470
rect 54392 27406 54444 27412
rect 56048 27464 56100 27470
rect 56048 27406 56100 27412
rect 54024 27328 54076 27334
rect 54024 27270 54076 27276
rect 54576 27328 54628 27334
rect 54576 27270 54628 27276
rect 56416 27328 56468 27334
rect 56416 27270 56468 27276
rect 54036 27062 54064 27270
rect 54024 27056 54076 27062
rect 54024 26998 54076 27004
rect 52644 26444 52696 26450
rect 52644 26386 52696 26392
rect 52460 26376 52512 26382
rect 52460 26318 52512 26324
rect 52920 26308 52972 26314
rect 52920 26250 52972 26256
rect 50632 25214 50752 25242
rect 50804 25288 50856 25294
rect 50804 25230 50856 25236
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50632 24750 50660 25214
rect 50712 25152 50764 25158
rect 50712 25094 50764 25100
rect 50620 24744 50672 24750
rect 50620 24686 50672 24692
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 49976 22636 50028 22642
rect 49976 22578 50028 22584
rect 49608 22432 49660 22438
rect 49608 22374 49660 22380
rect 49620 22098 49648 22374
rect 49608 22092 49660 22098
rect 49608 22034 49660 22040
rect 49988 20466 50016 22578
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 49976 20460 50028 20466
rect 49976 20402 50028 20408
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 50724 2650 50752 25094
rect 50988 20392 51040 20398
rect 50988 20334 51040 20340
rect 51000 3534 51028 20334
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 52932 2650 52960 26250
rect 54588 2650 54616 27270
rect 56428 2650 56456 27270
rect 58360 2650 58388 30126
rect 58716 30048 58768 30054
rect 58716 29990 58768 29996
rect 58728 29714 58756 29990
rect 60476 29850 60504 30126
rect 60464 29844 60516 29850
rect 60464 29786 60516 29792
rect 58716 29708 58768 29714
rect 58716 29650 58768 29656
rect 60660 29578 60688 37062
rect 61948 31482 61976 37062
rect 63040 31816 63092 31822
rect 63040 31758 63092 31764
rect 63500 31816 63552 31822
rect 63500 31758 63552 31764
rect 61936 31476 61988 31482
rect 61936 31418 61988 31424
rect 63052 31278 63080 31758
rect 63512 31482 63540 31758
rect 63880 31482 63908 37062
rect 65654 36476 65962 36496
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36400 65962 36420
rect 65654 35388 65962 35408
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35312 65962 35332
rect 65654 34300 65962 34320
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34224 65962 34244
rect 65654 33212 65962 33232
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33136 65962 33156
rect 65984 32428 66036 32434
rect 65984 32370 66036 32376
rect 65654 32124 65962 32144
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32048 65962 32068
rect 65996 32026 66024 32370
rect 65984 32020 66036 32026
rect 65984 31962 66036 31968
rect 66180 31754 66208 37062
rect 68204 33998 68232 37062
rect 69584 34746 69612 37062
rect 71516 35834 71544 37062
rect 73724 36922 73752 37062
rect 74736 36922 74764 37130
rect 75092 37120 75144 37126
rect 75092 37062 75144 37068
rect 75104 36922 75132 37062
rect 76760 36922 76788 39471
rect 77114 39200 77170 40000
rect 79046 39200 79102 40000
rect 76932 37256 76984 37262
rect 76932 37198 76984 37204
rect 73712 36916 73764 36922
rect 73712 36858 73764 36864
rect 74724 36916 74776 36922
rect 74724 36858 74776 36864
rect 75092 36916 75144 36922
rect 75092 36858 75144 36864
rect 76748 36916 76800 36922
rect 76748 36858 76800 36864
rect 76196 36780 76248 36786
rect 76196 36722 76248 36728
rect 73620 36712 73672 36718
rect 73620 36654 73672 36660
rect 73988 36712 74040 36718
rect 73988 36654 74040 36660
rect 75184 36712 75236 36718
rect 75184 36654 75236 36660
rect 73160 36100 73212 36106
rect 73160 36042 73212 36048
rect 73172 35834 73200 36042
rect 71504 35828 71556 35834
rect 71504 35770 71556 35776
rect 73160 35828 73212 35834
rect 73160 35770 73212 35776
rect 73252 35760 73304 35766
rect 73252 35702 73304 35708
rect 71412 35624 71464 35630
rect 71412 35566 71464 35572
rect 69572 34740 69624 34746
rect 69572 34682 69624 34688
rect 69848 34604 69900 34610
rect 69848 34546 69900 34552
rect 68376 34468 68428 34474
rect 68376 34410 68428 34416
rect 68388 34066 68416 34410
rect 68376 34060 68428 34066
rect 68376 34002 68428 34008
rect 68192 33992 68244 33998
rect 68192 33934 68244 33940
rect 67732 33856 67784 33862
rect 67732 33798 67784 33804
rect 68376 33856 68428 33862
rect 68376 33798 68428 33804
rect 67744 33522 67772 33798
rect 67732 33516 67784 33522
rect 67732 33458 67784 33464
rect 66168 31748 66220 31754
rect 66168 31690 66220 31696
rect 66076 31680 66128 31686
rect 66076 31622 66128 31628
rect 63500 31476 63552 31482
rect 63500 31418 63552 31424
rect 63868 31476 63920 31482
rect 63868 31418 63920 31424
rect 64144 31340 64196 31346
rect 64144 31282 64196 31288
rect 61844 31272 61896 31278
rect 61844 31214 61896 31220
rect 63040 31272 63092 31278
rect 63040 31214 63092 31220
rect 61016 31204 61068 31210
rect 61016 31146 61068 31152
rect 61028 30122 61056 31146
rect 61016 30116 61068 30122
rect 61016 30058 61068 30064
rect 61028 29714 61056 30058
rect 61016 29708 61068 29714
rect 61016 29650 61068 29656
rect 60648 29572 60700 29578
rect 60648 29514 60700 29520
rect 60740 29504 60792 29510
rect 60740 29446 60792 29452
rect 46664 2644 46716 2650
rect 46664 2586 46716 2592
rect 49148 2644 49200 2650
rect 49148 2586 49200 2592
rect 50712 2644 50764 2650
rect 50712 2586 50764 2592
rect 52920 2644 52972 2650
rect 52920 2586 52972 2592
rect 54576 2644 54628 2650
rect 54576 2586 54628 2592
rect 56416 2644 56468 2650
rect 56416 2586 56468 2592
rect 58348 2644 58400 2650
rect 58348 2586 58400 2592
rect 60752 2446 60780 29446
rect 61856 2650 61884 31214
rect 62120 31136 62172 31142
rect 62120 31078 62172 31084
rect 62132 30802 62160 31078
rect 62120 30796 62172 30802
rect 62120 30738 62172 30744
rect 64156 2650 64184 31282
rect 65654 31036 65962 31056
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30960 65962 30980
rect 65654 29948 65962 29968
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29872 65962 29892
rect 65654 28860 65962 28880
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28784 65962 28804
rect 65654 27772 65962 27792
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27696 65962 27716
rect 65654 26684 65962 26704
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26608 65962 26628
rect 65654 25596 65962 25616
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25520 65962 25540
rect 65654 24508 65962 24528
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24432 65962 24452
rect 65654 23420 65962 23440
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23344 65962 23364
rect 65654 22332 65962 22352
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22256 65962 22276
rect 65654 21244 65962 21264
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21168 65962 21188
rect 65654 20156 65962 20176
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20080 65962 20100
rect 65654 19068 65962 19088
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 18992 65962 19012
rect 65654 17980 65962 18000
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17904 65962 17924
rect 65654 16892 65962 16912
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16816 65962 16836
rect 65654 15804 65962 15824
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15728 65962 15748
rect 65654 14716 65962 14736
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14640 65962 14660
rect 65654 13628 65962 13648
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13552 65962 13572
rect 65654 12540 65962 12560
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12464 65962 12484
rect 65654 11452 65962 11472
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11376 65962 11396
rect 65654 10364 65962 10384
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10288 65962 10308
rect 65654 9276 65962 9296
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9200 65962 9220
rect 65654 8188 65962 8208
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8112 65962 8132
rect 65654 7100 65962 7120
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7024 65962 7044
rect 65654 6012 65962 6032
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5936 65962 5956
rect 65654 4924 65962 4944
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4848 65962 4868
rect 65654 3836 65962 3856
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3760 65962 3780
rect 65654 2748 65962 2768
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2672 65962 2692
rect 66088 2650 66116 31622
rect 68388 2650 68416 33798
rect 68928 33516 68980 33522
rect 68928 33458 68980 33464
rect 68940 31958 68968 33458
rect 68928 31952 68980 31958
rect 68928 31894 68980 31900
rect 69860 2650 69888 34546
rect 71424 2650 71452 35566
rect 73264 34474 73292 35702
rect 73252 34468 73304 34474
rect 73252 34410 73304 34416
rect 73264 33658 73292 34410
rect 73252 33652 73304 33658
rect 73252 33594 73304 33600
rect 73632 2650 73660 36654
rect 73804 36576 73856 36582
rect 73804 36518 73856 36524
rect 73816 36174 73844 36518
rect 73804 36168 73856 36174
rect 73804 36110 73856 36116
rect 74000 35766 74028 36654
rect 73988 35760 74040 35766
rect 73988 35702 74040 35708
rect 75196 2650 75224 36654
rect 76208 34202 76236 36722
rect 76748 36032 76800 36038
rect 76748 35974 76800 35980
rect 76196 34196 76248 34202
rect 76196 34138 76248 34144
rect 76760 33862 76788 35974
rect 76944 34746 76972 37198
rect 77128 36174 77156 39200
rect 77206 38584 77262 38593
rect 77206 38519 77262 38528
rect 77220 37466 77248 38519
rect 77850 37632 77906 37641
rect 77850 37567 77906 37576
rect 77864 37466 77892 37567
rect 77208 37460 77260 37466
rect 77208 37402 77260 37408
rect 77852 37460 77904 37466
rect 77852 37402 77904 37408
rect 77668 36780 77720 36786
rect 77668 36722 77720 36728
rect 77680 36242 77708 36722
rect 77850 36680 77906 36689
rect 77850 36615 77852 36624
rect 77904 36615 77906 36624
rect 77852 36586 77904 36592
rect 77668 36236 77720 36242
rect 77668 36178 77720 36184
rect 77116 36168 77168 36174
rect 77116 36110 77168 36116
rect 78036 36032 78088 36038
rect 78036 35974 78088 35980
rect 78048 35737 78076 35974
rect 78034 35728 78090 35737
rect 79060 35698 79088 39200
rect 78034 35663 78090 35672
rect 79048 35692 79100 35698
rect 79048 35634 79100 35640
rect 77760 35488 77812 35494
rect 77760 35430 77812 35436
rect 76932 34740 76984 34746
rect 76932 34682 76984 34688
rect 77208 34604 77260 34610
rect 77208 34546 77260 34552
rect 77300 34604 77352 34610
rect 77300 34546 77352 34552
rect 77220 34202 77248 34546
rect 77208 34196 77260 34202
rect 77208 34138 77260 34144
rect 77116 34060 77168 34066
rect 77116 34002 77168 34008
rect 76932 33924 76984 33930
rect 76932 33866 76984 33872
rect 76748 33856 76800 33862
rect 76748 33798 76800 33804
rect 76196 32904 76248 32910
rect 76196 32846 76248 32852
rect 76208 32230 76236 32846
rect 76196 32224 76248 32230
rect 76196 32166 76248 32172
rect 76196 27464 76248 27470
rect 76196 27406 76248 27412
rect 76208 26790 76236 27406
rect 76196 26784 76248 26790
rect 76196 26726 76248 26732
rect 76288 3392 76340 3398
rect 76288 3334 76340 3340
rect 76300 3194 76328 3334
rect 76944 3194 76972 33866
rect 77128 33386 77156 34002
rect 77208 33992 77260 33998
rect 77208 33934 77260 33940
rect 77220 33658 77248 33934
rect 77208 33652 77260 33658
rect 77208 33594 77260 33600
rect 77312 33454 77340 34546
rect 77772 33658 77800 35430
rect 77852 35080 77904 35086
rect 77852 35022 77904 35028
rect 77864 34678 77892 35022
rect 78036 34944 78088 34950
rect 78036 34886 78088 34892
rect 78048 34785 78076 34886
rect 78034 34776 78090 34785
rect 78034 34711 78090 34720
rect 77852 34672 77904 34678
rect 77852 34614 77904 34620
rect 77852 34400 77904 34406
rect 77852 34342 77904 34348
rect 77864 33969 77892 34342
rect 77850 33960 77906 33969
rect 77850 33895 77906 33904
rect 77760 33652 77812 33658
rect 77760 33594 77812 33600
rect 77944 33584 77996 33590
rect 77944 33526 77996 33532
rect 77300 33448 77352 33454
rect 77300 33390 77352 33396
rect 77116 33380 77168 33386
rect 77116 33322 77168 33328
rect 77128 20398 77156 33322
rect 77668 32428 77720 32434
rect 77668 32370 77720 32376
rect 77680 31822 77708 32370
rect 77852 32224 77904 32230
rect 77852 32166 77904 32172
rect 77864 32065 77892 32166
rect 77850 32056 77906 32065
rect 77850 31991 77906 32000
rect 77668 31816 77720 31822
rect 77668 31758 77720 31764
rect 77668 31340 77720 31346
rect 77668 31282 77720 31288
rect 77680 30734 77708 31282
rect 77852 31136 77904 31142
rect 77850 31104 77852 31113
rect 77904 31104 77906 31113
rect 77850 31039 77906 31048
rect 77668 30728 77720 30734
rect 77668 30670 77720 30676
rect 77850 30152 77906 30161
rect 77850 30087 77852 30096
rect 77904 30087 77906 30096
rect 77852 30058 77904 30064
rect 77852 28552 77904 28558
rect 77852 28494 77904 28500
rect 77864 27878 77892 28494
rect 77852 27872 77904 27878
rect 77852 27814 77904 27820
rect 77668 26988 77720 26994
rect 77668 26930 77720 26936
rect 77680 26314 77708 26930
rect 77852 26784 77904 26790
rect 77852 26726 77904 26732
rect 77864 26489 77892 26726
rect 77850 26480 77906 26489
rect 77850 26415 77906 26424
rect 77668 26308 77720 26314
rect 77668 26250 77720 26256
rect 77668 25900 77720 25906
rect 77668 25842 77720 25848
rect 77680 25158 77708 25842
rect 77852 25696 77904 25702
rect 77852 25638 77904 25644
rect 77864 25537 77892 25638
rect 77850 25528 77906 25537
rect 77850 25463 77906 25472
rect 77668 25152 77720 25158
rect 77668 25094 77720 25100
rect 77668 24812 77720 24818
rect 77668 24754 77720 24760
rect 77680 24070 77708 24754
rect 77852 24608 77904 24614
rect 77850 24576 77852 24585
rect 77904 24576 77906 24585
rect 77850 24511 77906 24520
rect 77668 24064 77720 24070
rect 77668 24006 77720 24012
rect 77850 23624 77906 23633
rect 77850 23559 77852 23568
rect 77904 23559 77906 23568
rect 77852 23530 77904 23536
rect 77484 22976 77536 22982
rect 77484 22918 77536 22924
rect 77496 22778 77524 22918
rect 77484 22772 77536 22778
rect 77484 22714 77536 22720
rect 77852 22024 77904 22030
rect 77852 21966 77904 21972
rect 77864 21690 77892 21966
rect 77852 21684 77904 21690
rect 77852 21626 77904 21632
rect 77116 20392 77168 20398
rect 77116 20334 77168 20340
rect 77852 20256 77904 20262
rect 77852 20198 77904 20204
rect 77864 19961 77892 20198
rect 77850 19952 77906 19961
rect 77850 19887 77906 19896
rect 77300 19372 77352 19378
rect 77300 19314 77352 19320
rect 77312 19174 77340 19314
rect 77300 19168 77352 19174
rect 77300 19110 77352 19116
rect 77852 19168 77904 19174
rect 77852 19110 77904 19116
rect 77312 18630 77340 19110
rect 77864 19009 77892 19110
rect 77850 19000 77906 19009
rect 77850 18935 77906 18944
rect 77300 18624 77352 18630
rect 77300 18566 77352 18572
rect 77852 18080 77904 18086
rect 77850 18048 77852 18057
rect 77904 18048 77906 18057
rect 77850 17983 77906 17992
rect 77852 17672 77904 17678
rect 77852 17614 77904 17620
rect 77864 16998 77892 17614
rect 77852 16992 77904 16998
rect 77852 16934 77904 16940
rect 77852 16584 77904 16590
rect 77852 16526 77904 16532
rect 77864 15910 77892 16526
rect 77852 15904 77904 15910
rect 77852 15846 77904 15852
rect 77852 13728 77904 13734
rect 77852 13670 77904 13676
rect 77864 13433 77892 13670
rect 77850 13424 77906 13433
rect 77850 13359 77906 13368
rect 77852 12640 77904 12646
rect 77852 12582 77904 12588
rect 77864 12481 77892 12582
rect 77850 12472 77906 12481
rect 77850 12407 77906 12416
rect 77850 11656 77906 11665
rect 77850 11591 77852 11600
rect 77904 11591 77906 11600
rect 77852 11562 77904 11568
rect 77956 10130 77984 33526
rect 78128 33516 78180 33522
rect 78128 33458 78180 33464
rect 78036 33040 78088 33046
rect 78034 33008 78036 33017
rect 78088 33008 78090 33017
rect 78034 32943 78090 32952
rect 78036 29504 78088 29510
rect 78036 29446 78088 29452
rect 78048 29209 78076 29446
rect 78034 29200 78090 29209
rect 78034 29135 78090 29144
rect 78036 28416 78088 28422
rect 78034 28384 78036 28393
rect 78088 28384 78090 28393
rect 78034 28319 78090 28328
rect 78034 27432 78090 27441
rect 78034 27367 78090 27376
rect 78048 27334 78076 27367
rect 78036 27328 78088 27334
rect 78036 27270 78088 27276
rect 78036 22976 78088 22982
rect 78036 22918 78088 22924
rect 78048 22817 78076 22918
rect 78034 22808 78090 22817
rect 78034 22743 78090 22752
rect 78036 21888 78088 21894
rect 78034 21856 78036 21865
rect 78088 21856 78090 21865
rect 78034 21791 78090 21800
rect 78034 20904 78090 20913
rect 78034 20839 78090 20848
rect 78048 20806 78076 20839
rect 78036 20800 78088 20806
rect 78036 20742 78088 20748
rect 78036 17536 78088 17542
rect 78036 17478 78088 17484
rect 78048 17241 78076 17478
rect 78034 17232 78090 17241
rect 78034 17167 78090 17176
rect 78036 16448 78088 16454
rect 78036 16390 78088 16396
rect 78048 16289 78076 16390
rect 78034 16280 78090 16289
rect 78034 16215 78090 16224
rect 78036 15360 78088 15366
rect 78034 15328 78036 15337
rect 78088 15328 78090 15337
rect 78034 15263 78090 15272
rect 78034 14376 78090 14385
rect 78034 14311 78090 14320
rect 78048 14278 78076 14311
rect 78036 14272 78088 14278
rect 78036 14214 78088 14220
rect 78036 11280 78088 11286
rect 78036 11222 78088 11228
rect 78048 10713 78076 11222
rect 78034 10704 78090 10713
rect 78034 10639 78090 10648
rect 77944 10124 77996 10130
rect 77944 10066 77996 10072
rect 77668 10056 77720 10062
rect 77668 9998 77720 10004
rect 77680 9761 77708 9998
rect 77666 9752 77722 9761
rect 77666 9687 77722 9696
rect 77668 8968 77720 8974
rect 77668 8910 77720 8916
rect 77576 8900 77628 8906
rect 77576 8842 77628 8848
rect 77208 7404 77260 7410
rect 77208 7346 77260 7352
rect 77220 6905 77248 7346
rect 77206 6896 77262 6905
rect 77206 6831 77262 6840
rect 77484 6316 77536 6322
rect 77484 6258 77536 6264
rect 77392 6248 77444 6254
rect 77392 6190 77444 6196
rect 77300 4548 77352 4554
rect 77300 4490 77352 4496
rect 77312 4146 77340 4490
rect 77300 4140 77352 4146
rect 77300 4082 77352 4088
rect 77404 3466 77432 6190
rect 77496 6089 77524 6258
rect 77482 6080 77538 6089
rect 77482 6015 77538 6024
rect 77484 5228 77536 5234
rect 77484 5170 77536 5176
rect 77496 5137 77524 5170
rect 77482 5128 77538 5137
rect 77482 5063 77538 5072
rect 77484 5024 77536 5030
rect 77484 4966 77536 4972
rect 77392 3460 77444 3466
rect 77392 3402 77444 3408
rect 76288 3188 76340 3194
rect 76288 3130 76340 3136
rect 76932 3188 76984 3194
rect 76932 3130 76984 3136
rect 77116 3052 77168 3058
rect 77116 2994 77168 3000
rect 77024 2984 77076 2990
rect 77024 2926 77076 2932
rect 61844 2644 61896 2650
rect 61844 2586 61896 2592
rect 64144 2644 64196 2650
rect 64144 2586 64196 2592
rect 66076 2644 66128 2650
rect 66076 2586 66128 2592
rect 68376 2644 68428 2650
rect 68376 2586 68428 2592
rect 69848 2644 69900 2650
rect 69848 2586 69900 2592
rect 71412 2644 71464 2650
rect 71412 2586 71464 2592
rect 73620 2644 73672 2650
rect 73620 2586 73672 2592
rect 75184 2644 75236 2650
rect 75184 2586 75236 2592
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 44732 2440 44784 2446
rect 44732 2382 44784 2388
rect 45284 2440 45336 2446
rect 45284 2382 45336 2388
rect 46664 2440 46716 2446
rect 46664 2382 46716 2388
rect 60740 2440 60792 2446
rect 60740 2382 60792 2388
rect 73344 2440 73396 2446
rect 73344 2382 73396 2388
rect 75184 2440 75236 2446
rect 75184 2382 75236 2388
rect 76564 2440 76616 2446
rect 76564 2382 76616 2388
rect 42812 800 42840 2382
rect 44744 800 44772 2382
rect 46676 800 46704 2382
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 50620 2372 50672 2378
rect 50620 2314 50672 2320
rect 52368 2372 52420 2378
rect 52368 2314 52420 2320
rect 54300 2372 54352 2378
rect 54300 2314 54352 2320
rect 56140 2372 56192 2378
rect 56140 2314 56192 2320
rect 58072 2372 58124 2378
rect 58072 2314 58124 2320
rect 60004 2372 60056 2378
rect 60004 2314 60056 2320
rect 61844 2372 61896 2378
rect 61844 2314 61896 2320
rect 63776 2372 63828 2378
rect 63776 2314 63828 2320
rect 65708 2372 65760 2378
rect 65708 2314 65760 2320
rect 67640 2372 67692 2378
rect 67640 2314 67692 2320
rect 69480 2372 69532 2378
rect 69480 2314 69532 2320
rect 71412 2372 71464 2378
rect 71412 2314 71464 2320
rect 48516 800 48544 2314
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50632 1170 50660 2314
rect 50448 1142 50660 1170
rect 50448 800 50476 1142
rect 52380 800 52408 2314
rect 54312 800 54340 2314
rect 56152 800 56180 2314
rect 58084 800 58112 2314
rect 60016 800 60044 2314
rect 61856 800 61884 2314
rect 63788 800 63816 2314
rect 65720 800 65748 2314
rect 67652 800 67680 2314
rect 69492 800 69520 2314
rect 71424 800 71452 2314
rect 73356 800 73384 2382
rect 75196 800 75224 2382
rect 938 0 994 800
rect 2778 0 2834 800
rect 4710 0 4766 800
rect 6642 0 6698 800
rect 8482 0 8538 800
rect 10414 0 10470 800
rect 12346 0 12402 800
rect 14278 0 14334 800
rect 16118 0 16174 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21822 0 21878 800
rect 23754 0 23810 800
rect 25686 0 25742 800
rect 27618 0 27674 800
rect 29458 0 29514 800
rect 31390 0 31446 800
rect 33322 0 33378 800
rect 35162 0 35218 800
rect 37094 0 37150 800
rect 39026 0 39082 800
rect 40958 0 41014 800
rect 42798 0 42854 800
rect 44730 0 44786 800
rect 46662 0 46718 800
rect 48502 0 48558 800
rect 50434 0 50490 800
rect 52366 0 52422 800
rect 54298 0 54354 800
rect 56138 0 56194 800
rect 58070 0 58126 800
rect 60002 0 60058 800
rect 61842 0 61898 800
rect 63774 0 63830 800
rect 65706 0 65762 800
rect 67638 0 67694 800
rect 69478 0 69534 800
rect 71410 0 71466 800
rect 73342 0 73398 800
rect 75182 0 75238 800
rect 76576 513 76604 2382
rect 77036 2281 77064 2926
rect 77022 2272 77078 2281
rect 77022 2207 77078 2216
rect 77128 800 77156 2994
rect 77208 2440 77260 2446
rect 77208 2382 77260 2388
rect 77220 1329 77248 2382
rect 77496 2038 77524 4966
rect 77588 2922 77616 8842
rect 77680 8809 77708 8910
rect 77666 8800 77722 8809
rect 77666 8735 77722 8744
rect 77668 7880 77720 7886
rect 77666 7848 77668 7857
rect 77720 7848 77722 7857
rect 77666 7783 77722 7792
rect 78036 7812 78088 7818
rect 78036 7754 78088 7760
rect 77852 7336 77904 7342
rect 77852 7278 77904 7284
rect 77668 4616 77720 4622
rect 77668 4558 77720 4564
rect 77680 4185 77708 4558
rect 77666 4176 77722 4185
rect 77666 4111 77722 4120
rect 77760 3596 77812 3602
rect 77760 3538 77812 3544
rect 77668 3528 77720 3534
rect 77668 3470 77720 3476
rect 77680 3233 77708 3470
rect 77666 3224 77722 3233
rect 77666 3159 77722 3168
rect 77772 3058 77800 3538
rect 77760 3052 77812 3058
rect 77760 2994 77812 3000
rect 77576 2916 77628 2922
rect 77576 2858 77628 2864
rect 77864 2582 77892 7278
rect 77944 3460 77996 3466
rect 77944 3402 77996 3408
rect 77956 3126 77984 3402
rect 78048 3398 78076 7754
rect 78140 4146 78168 33458
rect 79048 4208 79100 4214
rect 79048 4150 79100 4156
rect 78128 4140 78180 4146
rect 78128 4082 78180 4088
rect 78036 3392 78088 3398
rect 78036 3334 78088 3340
rect 77944 3120 77996 3126
rect 77944 3062 77996 3068
rect 77852 2576 77904 2582
rect 77852 2518 77904 2524
rect 77760 2372 77812 2378
rect 77760 2314 77812 2320
rect 77484 2032 77536 2038
rect 77484 1974 77536 1980
rect 77772 1970 77800 2314
rect 77760 1964 77812 1970
rect 77760 1906 77812 1912
rect 77206 1320 77262 1329
rect 77206 1255 77262 1264
rect 79060 800 79088 4150
rect 76562 504 76618 513
rect 76562 439 76618 448
rect 77114 0 77170 800
rect 79046 0 79102 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 76746 39480 76802 39536
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 77206 38528 77262 38584
rect 77850 37576 77906 37632
rect 77850 36644 77906 36680
rect 77850 36624 77852 36644
rect 77852 36624 77904 36644
rect 77904 36624 77906 36644
rect 78034 35672 78090 35728
rect 78034 34720 78090 34776
rect 77850 33904 77906 33960
rect 77850 32000 77906 32056
rect 77850 31084 77852 31104
rect 77852 31084 77904 31104
rect 77904 31084 77906 31104
rect 77850 31048 77906 31084
rect 77850 30116 77906 30152
rect 77850 30096 77852 30116
rect 77852 30096 77904 30116
rect 77904 30096 77906 30116
rect 77850 26424 77906 26480
rect 77850 25472 77906 25528
rect 77850 24556 77852 24576
rect 77852 24556 77904 24576
rect 77904 24556 77906 24576
rect 77850 24520 77906 24556
rect 77850 23588 77906 23624
rect 77850 23568 77852 23588
rect 77852 23568 77904 23588
rect 77904 23568 77906 23588
rect 77850 19896 77906 19952
rect 77850 18944 77906 19000
rect 77850 18028 77852 18048
rect 77852 18028 77904 18048
rect 77904 18028 77906 18048
rect 77850 17992 77906 18028
rect 77850 13368 77906 13424
rect 77850 12416 77906 12472
rect 77850 11620 77906 11656
rect 77850 11600 77852 11620
rect 77852 11600 77904 11620
rect 77904 11600 77906 11620
rect 78034 32988 78036 33008
rect 78036 32988 78088 33008
rect 78088 32988 78090 33008
rect 78034 32952 78090 32988
rect 78034 29144 78090 29200
rect 78034 28364 78036 28384
rect 78036 28364 78088 28384
rect 78088 28364 78090 28384
rect 78034 28328 78090 28364
rect 78034 27376 78090 27432
rect 78034 22752 78090 22808
rect 78034 21836 78036 21856
rect 78036 21836 78088 21856
rect 78088 21836 78090 21856
rect 78034 21800 78090 21836
rect 78034 20848 78090 20904
rect 78034 17176 78090 17232
rect 78034 16224 78090 16280
rect 78034 15308 78036 15328
rect 78036 15308 78088 15328
rect 78088 15308 78090 15328
rect 78034 15272 78090 15308
rect 78034 14320 78090 14376
rect 78034 10648 78090 10704
rect 77666 9696 77722 9752
rect 77206 6840 77262 6896
rect 77482 6024 77538 6080
rect 77482 5072 77538 5128
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 77022 2216 77078 2272
rect 77666 8744 77722 8800
rect 77666 7828 77668 7848
rect 77668 7828 77720 7848
rect 77720 7828 77722 7848
rect 77666 7792 77722 7828
rect 77666 4120 77722 4176
rect 77666 3168 77722 3224
rect 77206 1264 77262 1320
rect 76562 448 76618 504
<< metal3 >>
rect 76741 39538 76807 39541
rect 79200 39538 80000 39568
rect 76741 39536 80000 39538
rect 76741 39480 76746 39536
rect 76802 39480 80000 39536
rect 76741 39478 80000 39480
rect 76741 39475 76807 39478
rect 79200 39448 80000 39478
rect 77201 38586 77267 38589
rect 79200 38586 80000 38616
rect 77201 38584 80000 38586
rect 77201 38528 77206 38584
rect 77262 38528 80000 38584
rect 77201 38526 80000 38528
rect 77201 38523 77267 38526
rect 79200 38496 80000 38526
rect 77845 37634 77911 37637
rect 79200 37634 80000 37664
rect 77845 37632 80000 37634
rect 77845 37576 77850 37632
rect 77906 37576 80000 37632
rect 77845 37574 80000 37576
rect 77845 37571 77911 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 65648 37568 65968 37569
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 79200 37544 80000 37574
rect 65648 37503 65968 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 77845 36682 77911 36685
rect 79200 36682 80000 36712
rect 77845 36680 80000 36682
rect 77845 36624 77850 36680
rect 77906 36624 80000 36680
rect 77845 36622 80000 36624
rect 77845 36619 77911 36622
rect 79200 36592 80000 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 65648 36480 65968 36481
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36415 65968 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 78029 35730 78095 35733
rect 79200 35730 80000 35760
rect 78029 35728 80000 35730
rect 78029 35672 78034 35728
rect 78090 35672 80000 35728
rect 78029 35670 80000 35672
rect 78029 35667 78095 35670
rect 79200 35640 80000 35670
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 65648 35392 65968 35393
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 35327 65968 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 78029 34778 78095 34781
rect 79200 34778 80000 34808
rect 78029 34776 80000 34778
rect 78029 34720 78034 34776
rect 78090 34720 80000 34776
rect 78029 34718 80000 34720
rect 78029 34715 78095 34718
rect 79200 34688 80000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 65648 34304 65968 34305
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 34239 65968 34240
rect 77845 33962 77911 33965
rect 79200 33962 80000 33992
rect 77845 33960 80000 33962
rect 77845 33904 77850 33960
rect 77906 33904 80000 33960
rect 77845 33902 80000 33904
rect 77845 33899 77911 33902
rect 79200 33872 80000 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 65648 33216 65968 33217
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 33151 65968 33152
rect 78029 33010 78095 33013
rect 79200 33010 80000 33040
rect 78029 33008 80000 33010
rect 78029 32952 78034 33008
rect 78090 32952 80000 33008
rect 78029 32950 80000 32952
rect 78029 32947 78095 32950
rect 79200 32920 80000 32950
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 65648 32128 65968 32129
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 32063 65968 32064
rect 77845 32058 77911 32061
rect 79200 32058 80000 32088
rect 77845 32056 80000 32058
rect 77845 32000 77850 32056
rect 77906 32000 80000 32056
rect 77845 31998 80000 32000
rect 77845 31995 77911 31998
rect 79200 31968 80000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 77845 31106 77911 31109
rect 79200 31106 80000 31136
rect 77845 31104 80000 31106
rect 77845 31048 77850 31104
rect 77906 31048 80000 31104
rect 77845 31046 80000 31048
rect 77845 31043 77911 31046
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 65648 31040 65968 31041
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 79200 31016 80000 31046
rect 65648 30975 65968 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 77845 30154 77911 30157
rect 79200 30154 80000 30184
rect 77845 30152 80000 30154
rect 77845 30096 77850 30152
rect 77906 30096 80000 30152
rect 77845 30094 80000 30096
rect 77845 30091 77911 30094
rect 79200 30064 80000 30094
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 65648 29952 65968 29953
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 29887 65968 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 78029 29202 78095 29205
rect 79200 29202 80000 29232
rect 78029 29200 80000 29202
rect 78029 29144 78034 29200
rect 78090 29144 80000 29200
rect 78029 29142 80000 29144
rect 78029 29139 78095 29142
rect 79200 29112 80000 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 65648 28864 65968 28865
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 28799 65968 28800
rect 78029 28386 78095 28389
rect 79200 28386 80000 28416
rect 78029 28384 80000 28386
rect 78029 28328 78034 28384
rect 78090 28328 80000 28384
rect 78029 28326 80000 28328
rect 78029 28323 78095 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 79200 28296 80000 28326
rect 50288 28255 50608 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 65648 27776 65968 27777
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 27711 65968 27712
rect 78029 27434 78095 27437
rect 79200 27434 80000 27464
rect 78029 27432 80000 27434
rect 78029 27376 78034 27432
rect 78090 27376 80000 27432
rect 78029 27374 80000 27376
rect 78029 27371 78095 27374
rect 79200 27344 80000 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 65648 26688 65968 26689
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 26623 65968 26624
rect 77845 26482 77911 26485
rect 79200 26482 80000 26512
rect 77845 26480 80000 26482
rect 77845 26424 77850 26480
rect 77906 26424 80000 26480
rect 77845 26422 80000 26424
rect 77845 26419 77911 26422
rect 79200 26392 80000 26422
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 65648 25600 65968 25601
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 25535 65968 25536
rect 77845 25530 77911 25533
rect 79200 25530 80000 25560
rect 77845 25528 80000 25530
rect 77845 25472 77850 25528
rect 77906 25472 80000 25528
rect 77845 25470 80000 25472
rect 77845 25467 77911 25470
rect 79200 25440 80000 25470
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 77845 24578 77911 24581
rect 79200 24578 80000 24608
rect 77845 24576 80000 24578
rect 77845 24520 77850 24576
rect 77906 24520 80000 24576
rect 77845 24518 80000 24520
rect 77845 24515 77911 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 65648 24512 65968 24513
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 79200 24488 80000 24518
rect 65648 24447 65968 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 77845 23626 77911 23629
rect 79200 23626 80000 23656
rect 77845 23624 80000 23626
rect 77845 23568 77850 23624
rect 77906 23568 80000 23624
rect 77845 23566 80000 23568
rect 77845 23563 77911 23566
rect 79200 23536 80000 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 65648 23424 65968 23425
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 23359 65968 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 78029 22810 78095 22813
rect 79200 22810 80000 22840
rect 78029 22808 80000 22810
rect 78029 22752 78034 22808
rect 78090 22752 80000 22808
rect 78029 22750 80000 22752
rect 78029 22747 78095 22750
rect 79200 22720 80000 22750
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 65648 22336 65968 22337
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 22271 65968 22272
rect 78029 21858 78095 21861
rect 79200 21858 80000 21888
rect 78029 21856 80000 21858
rect 78029 21800 78034 21856
rect 78090 21800 80000 21856
rect 78029 21798 80000 21800
rect 78029 21795 78095 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 79200 21768 80000 21798
rect 50288 21727 50608 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 65648 21248 65968 21249
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 21183 65968 21184
rect 78029 20906 78095 20909
rect 79200 20906 80000 20936
rect 78029 20904 80000 20906
rect 78029 20848 78034 20904
rect 78090 20848 80000 20904
rect 78029 20846 80000 20848
rect 78029 20843 78095 20846
rect 79200 20816 80000 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 65648 20160 65968 20161
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 20095 65968 20096
rect 77845 19954 77911 19957
rect 79200 19954 80000 19984
rect 77845 19952 80000 19954
rect 77845 19896 77850 19952
rect 77906 19896 80000 19952
rect 77845 19894 80000 19896
rect 77845 19891 77911 19894
rect 79200 19864 80000 19894
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 65648 19072 65968 19073
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 19007 65968 19008
rect 77845 19002 77911 19005
rect 79200 19002 80000 19032
rect 77845 19000 80000 19002
rect 77845 18944 77850 19000
rect 77906 18944 80000 19000
rect 77845 18942 80000 18944
rect 77845 18939 77911 18942
rect 79200 18912 80000 18942
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 77845 18050 77911 18053
rect 79200 18050 80000 18080
rect 77845 18048 80000 18050
rect 77845 17992 77850 18048
rect 77906 17992 80000 18048
rect 77845 17990 80000 17992
rect 77845 17987 77911 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 65648 17984 65968 17985
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 79200 17960 80000 17990
rect 65648 17919 65968 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 78029 17234 78095 17237
rect 79200 17234 80000 17264
rect 78029 17232 80000 17234
rect 78029 17176 78034 17232
rect 78090 17176 80000 17232
rect 78029 17174 80000 17176
rect 78029 17171 78095 17174
rect 79200 17144 80000 17174
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 65648 16896 65968 16897
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 16831 65968 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 78029 16282 78095 16285
rect 79200 16282 80000 16312
rect 78029 16280 80000 16282
rect 78029 16224 78034 16280
rect 78090 16224 80000 16280
rect 78029 16222 80000 16224
rect 78029 16219 78095 16222
rect 79200 16192 80000 16222
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 65648 15808 65968 15809
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 15743 65968 15744
rect 78029 15330 78095 15333
rect 79200 15330 80000 15360
rect 78029 15328 80000 15330
rect 78029 15272 78034 15328
rect 78090 15272 80000 15328
rect 78029 15270 80000 15272
rect 78029 15267 78095 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 79200 15240 80000 15270
rect 50288 15199 50608 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 65648 14720 65968 14721
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 14655 65968 14656
rect 78029 14378 78095 14381
rect 79200 14378 80000 14408
rect 78029 14376 80000 14378
rect 78029 14320 78034 14376
rect 78090 14320 80000 14376
rect 78029 14318 80000 14320
rect 78029 14315 78095 14318
rect 79200 14288 80000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 65648 13632 65968 13633
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 13567 65968 13568
rect 77845 13426 77911 13429
rect 79200 13426 80000 13456
rect 77845 13424 80000 13426
rect 77845 13368 77850 13424
rect 77906 13368 80000 13424
rect 77845 13366 80000 13368
rect 77845 13363 77911 13366
rect 79200 13336 80000 13366
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 65648 12544 65968 12545
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 12479 65968 12480
rect 77845 12474 77911 12477
rect 79200 12474 80000 12504
rect 77845 12472 80000 12474
rect 77845 12416 77850 12472
rect 77906 12416 80000 12472
rect 77845 12414 80000 12416
rect 77845 12411 77911 12414
rect 79200 12384 80000 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 77845 11658 77911 11661
rect 79200 11658 80000 11688
rect 77845 11656 80000 11658
rect 77845 11600 77850 11656
rect 77906 11600 80000 11656
rect 77845 11598 80000 11600
rect 77845 11595 77911 11598
rect 79200 11568 80000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 65648 11456 65968 11457
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 11391 65968 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 78029 10706 78095 10709
rect 79200 10706 80000 10736
rect 78029 10704 80000 10706
rect 78029 10648 78034 10704
rect 78090 10648 80000 10704
rect 78029 10646 80000 10648
rect 78029 10643 78095 10646
rect 79200 10616 80000 10646
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 65648 10368 65968 10369
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 10303 65968 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 77661 9754 77727 9757
rect 79200 9754 80000 9784
rect 77661 9752 80000 9754
rect 77661 9696 77666 9752
rect 77722 9696 80000 9752
rect 77661 9694 80000 9696
rect 77661 9691 77727 9694
rect 79200 9664 80000 9694
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 65648 9280 65968 9281
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 9215 65968 9216
rect 77661 8802 77727 8805
rect 79200 8802 80000 8832
rect 77661 8800 80000 8802
rect 77661 8744 77666 8800
rect 77722 8744 80000 8800
rect 77661 8742 80000 8744
rect 77661 8739 77727 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 79200 8712 80000 8742
rect 50288 8671 50608 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 65648 8192 65968 8193
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 8127 65968 8128
rect 77661 7850 77727 7853
rect 79200 7850 80000 7880
rect 77661 7848 80000 7850
rect 77661 7792 77666 7848
rect 77722 7792 80000 7848
rect 77661 7790 80000 7792
rect 77661 7787 77727 7790
rect 79200 7760 80000 7790
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 65648 7104 65968 7105
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 7039 65968 7040
rect 77201 6898 77267 6901
rect 79200 6898 80000 6928
rect 77201 6896 80000 6898
rect 77201 6840 77206 6896
rect 77262 6840 80000 6896
rect 77201 6838 80000 6840
rect 77201 6835 77267 6838
rect 79200 6808 80000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 77477 6082 77543 6085
rect 79200 6082 80000 6112
rect 77477 6080 80000 6082
rect 77477 6024 77482 6080
rect 77538 6024 80000 6080
rect 77477 6022 80000 6024
rect 77477 6019 77543 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 65648 6016 65968 6017
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 79200 5992 80000 6022
rect 65648 5951 65968 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 77477 5130 77543 5133
rect 79200 5130 80000 5160
rect 77477 5128 80000 5130
rect 77477 5072 77482 5128
rect 77538 5072 80000 5128
rect 77477 5070 80000 5072
rect 77477 5067 77543 5070
rect 79200 5040 80000 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 65648 4928 65968 4929
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 4863 65968 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 77661 4178 77727 4181
rect 79200 4178 80000 4208
rect 77661 4176 80000 4178
rect 77661 4120 77666 4176
rect 77722 4120 80000 4176
rect 77661 4118 80000 4120
rect 77661 4115 77727 4118
rect 79200 4088 80000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 65648 3840 65968 3841
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 3775 65968 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 77661 3226 77727 3229
rect 79200 3226 80000 3256
rect 77661 3224 80000 3226
rect 77661 3168 77666 3224
rect 77722 3168 80000 3224
rect 77661 3166 80000 3168
rect 77661 3163 77727 3166
rect 79200 3136 80000 3166
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 65648 2752 65968 2753
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2687 65968 2688
rect 77017 2274 77083 2277
rect 79200 2274 80000 2304
rect 77017 2272 80000 2274
rect 77017 2216 77022 2272
rect 77078 2216 80000 2272
rect 77017 2214 80000 2216
rect 77017 2211 77083 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 79200 2184 80000 2214
rect 50288 2143 50608 2144
rect 77201 1322 77267 1325
rect 79200 1322 80000 1352
rect 77201 1320 80000 1322
rect 77201 1264 77206 1320
rect 77262 1264 80000 1320
rect 77201 1262 80000 1264
rect 77201 1259 77267 1262
rect 79200 1232 80000 1262
rect 76557 506 76623 509
rect 79200 506 80000 536
rect 76557 504 80000 506
rect 76557 448 76562 504
rect 76618 448 80000 504
rect 76557 446 80000 448
rect 76557 443 76623 446
rect 79200 416 80000 446
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 37024 50608 37584
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 37568 65968 37584
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 77464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 77280 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 77280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 77280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 77280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 77280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform -1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform -1 0 14168 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform -1 0 15088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform -1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform 1 0 77464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122
timestamp 1644511149
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_127
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 1644511149
transform 1 0 14720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_256
timestamp 1644511149
transform 1 0 24656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1644511149
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_292
timestamp 1644511149
transform 1 0 27968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_312
timestamp 1644511149
transform 1 0 29808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_324
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_340
timestamp 1644511149
transform 1 0 32384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_348
timestamp 1644511149
transform 1 0 33120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_381
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1644511149
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1644511149
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_431
timestamp 1644511149
transform 1 0 40756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1644511149
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1644511149
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_453
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_464
timestamp 1644511149
transform 1 0 43792 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_487
timestamp 1644511149
transform 1 0 45908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_499
timestamp 1644511149
transform 1 0 47012 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1644511149
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1644511149
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1644511149
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1644511149
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_541
timestamp 1644511149
transform 1 0 50876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1644511149
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1644511149
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_565
timestamp 1644511149
transform 1 0 53084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_577
timestamp 1644511149
transform 1 0 54188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_583
timestamp 1644511149
transform 1 0 54740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1644511149
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_597
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_603
timestamp 1644511149
transform 1 0 56580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1644511149
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_624
timestamp 1644511149
transform 1 0 58512 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_636
timestamp 1644511149
transform 1 0 59616 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_649
timestamp 1644511149
transform 1 0 60812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_665
timestamp 1644511149
transform 1 0 62284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1644511149
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_673
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_681
timestamp 1644511149
transform 1 0 63756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_686
timestamp 1644511149
transform 1 0 64216 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_698
timestamp 1644511149
transform 1 0 65320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_701
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_707
timestamp 1644511149
transform 1 0 66148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_719
timestamp 1644511149
transform 1 0 67252 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 1644511149
transform 1 0 67988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_733
timestamp 1644511149
transform 1 0 68540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_741
timestamp 1644511149
transform 1 0 69276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_748
timestamp 1644511149
transform 1 0 69920 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_757
timestamp 1644511149
transform 1 0 70748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_769
timestamp 1644511149
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1644511149
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_785
timestamp 1644511149
transform 1 0 73324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_790
timestamp 1644511149
transform 1 0 73784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_802
timestamp 1644511149
transform 1 0 74888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 1644511149
transform 1 0 75440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_813
timestamp 1644511149
transform 1 0 75900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_819
timestamp 1644511149
transform 1 0 76452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_826
timestamp 1644511149
transform 1 0 77096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_836
timestamp 1644511149
transform 1 0 78016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_841
timestamp 1644511149
transform 1 0 78476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1644511149
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1644511149
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_158
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1644511149
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1644511149
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1644511149
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1644511149
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_433
timestamp 1644511149
transform 1 0 40940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1644511149
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_641
timestamp 1644511149
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1644511149
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1644511149
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1644511149
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1644511149
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_697
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_709
timestamp 1644511149
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1644511149
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1644511149
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_729
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_741
timestamp 1644511149
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_753
timestamp 1644511149
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_765
timestamp 1644511149
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1644511149
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1644511149
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_785
timestamp 1644511149
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_797
timestamp 1644511149
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_809
timestamp 1644511149
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_821
timestamp 1644511149
transform 1 0 76636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_826
timestamp 1644511149
transform 1 0 77096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_836
timestamp 1644511149
transform 1 0 78016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_841
timestamp 1644511149
transform 1 0 78476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1644511149
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1644511149
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1644511149
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1644511149
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1644511149
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_681
timestamp 1644511149
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1644511149
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1644511149
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_713
timestamp 1644511149
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_725
timestamp 1644511149
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_737
timestamp 1644511149
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1644511149
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1644511149
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_757
timestamp 1644511149
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_769
timestamp 1644511149
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_781
timestamp 1644511149
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_793
timestamp 1644511149
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1644511149
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1644511149
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_813
timestamp 1644511149
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_825
timestamp 1644511149
transform 1 0 77004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_831
timestamp 1644511149
transform 1 0 77556 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_838
timestamp 1644511149
transform 1 0 78200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_653
timestamp 1644511149
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1644511149
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1644511149
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_673
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_685
timestamp 1644511149
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_697
timestamp 1644511149
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_709
timestamp 1644511149
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1644511149
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1644511149
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_729
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_741
timestamp 1644511149
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_753
timestamp 1644511149
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_765
timestamp 1644511149
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1644511149
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1644511149
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_785
timestamp 1644511149
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_797
timestamp 1644511149
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_809
timestamp 1644511149
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_821
timestamp 1644511149
transform 1 0 76636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_829
timestamp 1644511149
transform 1 0 77372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_836
timestamp 1644511149
transform 1 0 78016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_841
timestamp 1644511149
transform 1 0 78476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_669
timestamp 1644511149
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_681
timestamp 1644511149
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1644511149
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1644511149
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_725
timestamp 1644511149
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_737
timestamp 1644511149
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1644511149
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1644511149
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_757
timestamp 1644511149
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_769
timestamp 1644511149
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_781
timestamp 1644511149
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_793
timestamp 1644511149
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1644511149
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1644511149
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_813
timestamp 1644511149
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_825
timestamp 1644511149
transform 1 0 77004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_831
timestamp 1644511149
transform 1 0 77556 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_838
timestamp 1644511149
transform 1 0 78200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_673
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1644511149
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_697
timestamp 1644511149
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_709
timestamp 1644511149
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1644511149
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1644511149
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_741
timestamp 1644511149
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_753
timestamp 1644511149
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_765
timestamp 1644511149
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1644511149
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1644511149
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_785
timestamp 1644511149
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_797
timestamp 1644511149
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_809
timestamp 1644511149
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_821
timestamp 1644511149
transform 1 0 76636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_829
timestamp 1644511149
transform 1 0 77372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_836
timestamp 1644511149
transform 1 0 78016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_841
timestamp 1644511149
transform 1 0 78476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_713
timestamp 1644511149
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_737
timestamp 1644511149
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1644511149
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1644511149
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_757
timestamp 1644511149
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_769
timestamp 1644511149
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_781
timestamp 1644511149
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_793
timestamp 1644511149
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1644511149
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1644511149
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_813
timestamp 1644511149
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_825
timestamp 1644511149
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_837
timestamp 1644511149
transform 1 0 78108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_841
timestamp 1644511149
transform 1 0 78476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1644511149
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1644511149
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1644511149
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_741
timestamp 1644511149
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_753
timestamp 1644511149
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_765
timestamp 1644511149
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1644511149
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1644511149
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_785
timestamp 1644511149
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_797
timestamp 1644511149
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_809
timestamp 1644511149
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_821
timestamp 1644511149
transform 1 0 76636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_829
timestamp 1644511149
transform 1 0 77372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_836
timestamp 1644511149
transform 1 0 78016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_841
timestamp 1644511149
transform 1 0 78476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_725
timestamp 1644511149
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_737
timestamp 1644511149
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1644511149
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1644511149
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_757
timestamp 1644511149
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_769
timestamp 1644511149
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1644511149
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_793
timestamp 1644511149
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1644511149
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1644511149
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_813
timestamp 1644511149
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_825
timestamp 1644511149
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_837
timestamp 1644511149
transform 1 0 78108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_841
timestamp 1644511149
transform 1 0 78476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1644511149
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_741
timestamp 1644511149
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_753
timestamp 1644511149
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_765
timestamp 1644511149
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1644511149
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1644511149
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_785
timestamp 1644511149
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_797
timestamp 1644511149
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_809
timestamp 1644511149
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_821
timestamp 1644511149
transform 1 0 76636 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_829
timestamp 1644511149
transform 1 0 77372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_836
timestamp 1644511149
transform 1 0 78016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_841
timestamp 1644511149
transform 1 0 78476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1644511149
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_101
timestamp 1644511149
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_113
timestamp 1644511149
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_125
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1644511149
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_725
timestamp 1644511149
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_737
timestamp 1644511149
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1644511149
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1644511149
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_757
timestamp 1644511149
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_769
timestamp 1644511149
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_781
timestamp 1644511149
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_793
timestamp 1644511149
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1644511149
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1644511149
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_813
timestamp 1644511149
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_825
timestamp 1644511149
transform 1 0 77004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_831
timestamp 1644511149
transform 1 0 77556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_838
timestamp 1644511149
transform 1 0 78200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1644511149
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_741
timestamp 1644511149
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_753
timestamp 1644511149
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_765
timestamp 1644511149
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1644511149
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1644511149
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_785
timestamp 1644511149
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_797
timestamp 1644511149
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_809
timestamp 1644511149
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_821
timestamp 1644511149
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1644511149
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1644511149
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_841
timestamp 1644511149
transform 1 0 78476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_73
timestamp 1644511149
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_89
timestamp 1644511149
transform 1 0 9292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_101
timestamp 1644511149
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_113
timestamp 1644511149
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1644511149
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_737
timestamp 1644511149
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1644511149
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1644511149
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_757
timestamp 1644511149
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_769
timestamp 1644511149
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_781
timestamp 1644511149
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_793
timestamp 1644511149
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1644511149
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1644511149
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_813
timestamp 1644511149
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_825
timestamp 1644511149
transform 1 0 77004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_831
timestamp 1644511149
transform 1 0 77556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_838
timestamp 1644511149
transform 1 0 78200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_741
timestamp 1644511149
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_753
timestamp 1644511149
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_765
timestamp 1644511149
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1644511149
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1644511149
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_785
timestamp 1644511149
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_797
timestamp 1644511149
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_809
timestamp 1644511149
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_821
timestamp 1644511149
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1644511149
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1644511149
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_841
timestamp 1644511149
transform 1 0 78476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_737
timestamp 1644511149
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1644511149
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1644511149
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_757
timestamp 1644511149
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_769
timestamp 1644511149
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_781
timestamp 1644511149
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_793
timestamp 1644511149
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1644511149
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1644511149
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_813
timestamp 1644511149
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_825
timestamp 1644511149
transform 1 0 77004 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_831
timestamp 1644511149
transform 1 0 77556 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_838
timestamp 1644511149
transform 1 0 78200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_741
timestamp 1644511149
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_753
timestamp 1644511149
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_765
timestamp 1644511149
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1644511149
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1644511149
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_785
timestamp 1644511149
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_797
timestamp 1644511149
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_809
timestamp 1644511149
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_821
timestamp 1644511149
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1644511149
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1644511149
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_841
timestamp 1644511149
transform 1 0 78476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1644511149
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_737
timestamp 1644511149
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1644511149
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1644511149
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_757
timestamp 1644511149
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_769
timestamp 1644511149
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_781
timestamp 1644511149
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_793
timestamp 1644511149
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1644511149
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1644511149
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_813
timestamp 1644511149
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_825
timestamp 1644511149
transform 1 0 77004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_833
timestamp 1644511149
transform 1 0 77740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_838
timestamp 1644511149
transform 1 0 78200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_234
timestamp 1644511149
transform 1 0 22632 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_252
timestamp 1644511149
transform 1 0 24288 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_264
timestamp 1644511149
transform 1 0 25392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_741
timestamp 1644511149
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_753
timestamp 1644511149
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_765
timestamp 1644511149
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1644511149
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1644511149
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_785
timestamp 1644511149
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_797
timestamp 1644511149
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_809
timestamp 1644511149
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_821
timestamp 1644511149
transform 1 0 76636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_829
timestamp 1644511149
transform 1 0 77372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_836
timestamp 1644511149
transform 1 0 78016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_841
timestamp 1644511149
transform 1 0 78476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_259
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_271
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_283
timestamp 1644511149
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_295
timestamp 1644511149
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_737
timestamp 1644511149
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1644511149
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1644511149
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_757
timestamp 1644511149
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_769
timestamp 1644511149
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_781
timestamp 1644511149
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_793
timestamp 1644511149
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1644511149
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1644511149
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_813
timestamp 1644511149
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_825
timestamp 1644511149
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_837
timestamp 1644511149
transform 1 0 78108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_841
timestamp 1644511149
transform 1 0 78476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_741
timestamp 1644511149
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_753
timestamp 1644511149
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_765
timestamp 1644511149
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1644511149
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1644511149
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_785
timestamp 1644511149
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_797
timestamp 1644511149
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_809
timestamp 1644511149
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_821
timestamp 1644511149
transform 1 0 76636 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_827
timestamp 1644511149
transform 1 0 77188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_830
timestamp 1644511149
transform 1 0 77464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1644511149
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_841
timestamp 1644511149
transform 1 0 78476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_283
timestamp 1644511149
transform 1 0 27140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_295
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_725
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_737
timestamp 1644511149
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1644511149
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1644511149
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_757
timestamp 1644511149
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_769
timestamp 1644511149
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_781
timestamp 1644511149
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_793
timestamp 1644511149
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1644511149
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1644511149
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_813
timestamp 1644511149
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_825
timestamp 1644511149
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_837
timestamp 1644511149
transform 1 0 78108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_841
timestamp 1644511149
transform 1 0 78476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1644511149
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_148
timestamp 1644511149
transform 1 0 14720 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_292
timestamp 1644511149
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_304
timestamp 1644511149
transform 1 0 29072 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_316
timestamp 1644511149
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_328
timestamp 1644511149
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_741
timestamp 1644511149
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_753
timestamp 1644511149
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_765
timestamp 1644511149
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1644511149
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1644511149
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_785
timestamp 1644511149
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_797
timestamp 1644511149
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_809
timestamp 1644511149
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_821
timestamp 1644511149
transform 1 0 76636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_827
timestamp 1644511149
transform 1 0 77188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_830
timestamp 1644511149
transform 1 0 77464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_836
timestamp 1644511149
transform 1 0 78016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_841
timestamp 1644511149
transform 1 0 78476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_148
timestamp 1644511149
transform 1 0 14720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_285
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_725
timestamp 1644511149
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_737
timestamp 1644511149
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1644511149
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1644511149
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_757
timestamp 1644511149
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_769
timestamp 1644511149
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_781
timestamp 1644511149
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_793
timestamp 1644511149
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1644511149
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1644511149
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_813
timestamp 1644511149
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_825
timestamp 1644511149
transform 1 0 77004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_833
timestamp 1644511149
transform 1 0 77740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_838
timestamp 1644511149
transform 1 0 78200 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_133
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp 1644511149
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_156
timestamp 1644511149
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_173
timestamp 1644511149
transform 1 0 17020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_185
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_190
timestamp 1644511149
transform 1 0 18584 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_673
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1644511149
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_697
timestamp 1644511149
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_709
timestamp 1644511149
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1644511149
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1644511149
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_741
timestamp 1644511149
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_753
timestamp 1644511149
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_765
timestamp 1644511149
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1644511149
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1644511149
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_785
timestamp 1644511149
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_797
timestamp 1644511149
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_809
timestamp 1644511149
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_821
timestamp 1644511149
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1644511149
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1644511149
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_841
timestamp 1644511149
transform 1 0 78476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_146
timestamp 1644511149
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_158
timestamp 1644511149
transform 1 0 15640 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_170
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_182
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1644511149
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_315
timestamp 1644511149
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_322
timestamp 1644511149
transform 1 0 30728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_334
timestamp 1644511149
transform 1 0 31832 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_346
timestamp 1644511149
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1644511149
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1644511149
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1644511149
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1644511149
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_737
timestamp 1644511149
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1644511149
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1644511149
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_757
timestamp 1644511149
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_769
timestamp 1644511149
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_781
timestamp 1644511149
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_793
timestamp 1644511149
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1644511149
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1644511149
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_813
timestamp 1644511149
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_825
timestamp 1644511149
transform 1 0 77004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_833
timestamp 1644511149
transform 1 0 77740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_838
timestamp 1644511149
transform 1 0 78200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1644511149
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1644511149
transform 1 0 32660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1644511149
transform 1 0 33764 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1644511149
transform 1 0 34868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1644511149
transform 1 0 35972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_741
timestamp 1644511149
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_753
timestamp 1644511149
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_765
timestamp 1644511149
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1644511149
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1644511149
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_785
timestamp 1644511149
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_797
timestamp 1644511149
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_809
timestamp 1644511149
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_821
timestamp 1644511149
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1644511149
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1644511149
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_841
timestamp 1644511149
transform 1 0 78476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_325
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_335
timestamp 1644511149
transform 1 0 31924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_347
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_737
timestamp 1644511149
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1644511149
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1644511149
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_757
timestamp 1644511149
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_769
timestamp 1644511149
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_781
timestamp 1644511149
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_793
timestamp 1644511149
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1644511149
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1644511149
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_813
timestamp 1644511149
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_825
timestamp 1644511149
transform 1 0 77004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_833
timestamp 1644511149
transform 1 0 77740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_838
timestamp 1644511149
transform 1 0 78200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_345
timestamp 1644511149
transform 1 0 32844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_356
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_364
timestamp 1644511149
transform 1 0 34592 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_376
timestamp 1644511149
transform 1 0 35696 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_641
timestamp 1644511149
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_653
timestamp 1644511149
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1644511149
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1644511149
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1644511149
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1644511149
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1644511149
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_741
timestamp 1644511149
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_753
timestamp 1644511149
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_765
timestamp 1644511149
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1644511149
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1644511149
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_785
timestamp 1644511149
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_797
timestamp 1644511149
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_809
timestamp 1644511149
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_821
timestamp 1644511149
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1644511149
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1644511149
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_841
timestamp 1644511149
transform 1 0 78476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_376
timestamp 1644511149
transform 1 0 35696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1644511149
transform 1 0 36432 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_396
timestamp 1644511149
transform 1 0 37536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_408
timestamp 1644511149
transform 1 0 38640 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_725
timestamp 1644511149
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_737
timestamp 1644511149
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1644511149
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1644511149
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_757
timestamp 1644511149
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_769
timestamp 1644511149
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_781
timestamp 1644511149
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_793
timestamp 1644511149
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1644511149
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1644511149
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_813
timestamp 1644511149
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_825
timestamp 1644511149
transform 1 0 77004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_833
timestamp 1644511149
transform 1 0 77740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_838
timestamp 1644511149
transform 1 0 78200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_402
timestamp 1644511149
transform 1 0 38088 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_414
timestamp 1644511149
transform 1 0 39192 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_426
timestamp 1644511149
transform 1 0 40296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_438
timestamp 1644511149
transform 1 0 41400 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1644511149
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_741
timestamp 1644511149
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_753
timestamp 1644511149
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_765
timestamp 1644511149
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1644511149
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1644511149
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_785
timestamp 1644511149
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_797
timestamp 1644511149
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_809
timestamp 1644511149
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_821
timestamp 1644511149
transform 1 0 76636 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_827
timestamp 1644511149
transform 1 0 77188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_830
timestamp 1644511149
transform 1 0 77464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_836
timestamp 1644511149
transform 1 0 78016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_841
timestamp 1644511149
transform 1 0 78476 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1644511149
transform 1 0 38640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_625
timestamp 1644511149
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1644511149
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1644511149
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_725
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_737
timestamp 1644511149
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1644511149
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1644511149
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_757
timestamp 1644511149
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_769
timestamp 1644511149
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_781
timestamp 1644511149
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_793
timestamp 1644511149
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1644511149
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1644511149
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_813
timestamp 1644511149
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_825
timestamp 1644511149
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_837
timestamp 1644511149
transform 1 0 78108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_841
timestamp 1644511149
transform 1 0 78476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1644511149
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1644511149
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1644511149
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1644511149
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_741
timestamp 1644511149
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_753
timestamp 1644511149
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_765
timestamp 1644511149
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1644511149
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1644511149
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_785
timestamp 1644511149
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_797
timestamp 1644511149
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_809
timestamp 1644511149
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_821
timestamp 1644511149
transform 1 0 76636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_827
timestamp 1644511149
transform 1 0 77188 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_830
timestamp 1644511149
transform 1 0 77464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_836
timestamp 1644511149
transform 1 0 78016 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_841
timestamp 1644511149
transform 1 0 78476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_681
timestamp 1644511149
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1644511149
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_737
timestamp 1644511149
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1644511149
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1644511149
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_757
timestamp 1644511149
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_769
timestamp 1644511149
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_781
timestamp 1644511149
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_793
timestamp 1644511149
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1644511149
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1644511149
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_813
timestamp 1644511149
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_825
timestamp 1644511149
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_837
timestamp 1644511149
transform 1 0 78108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_841
timestamp 1644511149
transform 1 0 78476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_423
timestamp 1644511149
transform 1 0 40020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_435
timestamp 1644511149
transform 1 0 41124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_440
timestamp 1644511149
transform 1 0 41584 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_547
timestamp 1644511149
transform 1 0 51428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1644511149
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_673
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_685
timestamp 1644511149
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_697
timestamp 1644511149
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_709
timestamp 1644511149
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1644511149
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1644511149
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_729
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_741
timestamp 1644511149
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_753
timestamp 1644511149
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_765
timestamp 1644511149
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1644511149
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1644511149
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_785
timestamp 1644511149
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_797
timestamp 1644511149
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_809
timestamp 1644511149
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_821
timestamp 1644511149
transform 1 0 76636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_829
timestamp 1644511149
transform 1 0 77372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_836
timestamp 1644511149
transform 1 0 78016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_841
timestamp 1644511149
transform 1 0 78476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_430
timestamp 1644511149
transform 1 0 40664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_443
timestamp 1644511149
transform 1 0 41860 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_455
timestamp 1644511149
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_467
timestamp 1644511149
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1644511149
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1644511149
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1644511149
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1644511149
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_737
timestamp 1644511149
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1644511149
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1644511149
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_757
timestamp 1644511149
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_769
timestamp 1644511149
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_781
timestamp 1644511149
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_793
timestamp 1644511149
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1644511149
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1644511149
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_813
timestamp 1644511149
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_825
timestamp 1644511149
transform 1 0 77004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_829
timestamp 1644511149
transform 1 0 77372 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_832
timestamp 1644511149
transform 1 0 77648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_838
timestamp 1644511149
transform 1 0 78200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1644511149
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1644511149
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_709
timestamp 1644511149
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1644511149
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1644511149
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_741
timestamp 1644511149
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_753
timestamp 1644511149
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_765
timestamp 1644511149
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1644511149
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1644511149
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_785
timestamp 1644511149
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_797
timestamp 1644511149
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_809
timestamp 1644511149
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_821
timestamp 1644511149
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1644511149
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1644511149
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_841
timestamp 1644511149
transform 1 0 78476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_428
timestamp 1644511149
transform 1 0 40480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_440
timestamp 1644511149
transform 1 0 41584 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_448
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_459
timestamp 1644511149
transform 1 0 43332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_467
timestamp 1644511149
transform 1 0 44068 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_481
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_493
timestamp 1644511149
transform 1 0 46460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_505
timestamp 1644511149
transform 1 0 47564 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_517
timestamp 1644511149
transform 1 0 48668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_529
timestamp 1644511149
transform 1 0 49772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_625
timestamp 1644511149
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1644511149
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1644511149
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1644511149
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1644511149
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1644511149
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1644511149
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_725
timestamp 1644511149
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_737
timestamp 1644511149
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1644511149
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1644511149
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_757
timestamp 1644511149
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_769
timestamp 1644511149
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_781
timestamp 1644511149
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_793
timestamp 1644511149
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1644511149
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1644511149
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_813
timestamp 1644511149
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_825
timestamp 1644511149
transform 1 0 77004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_833
timestamp 1644511149
transform 1 0 77740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_838
timestamp 1644511149
transform 1 0 78200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_469
timestamp 1644511149
transform 1 0 44252 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_480
timestamp 1644511149
transform 1 0 45264 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_488
timestamp 1644511149
transform 1 0 46000 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_499
timestamp 1644511149
transform 1 0 47012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_536
timestamp 1644511149
transform 1 0 50416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_548
timestamp 1644511149
transform 1 0 51520 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1644511149
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_741
timestamp 1644511149
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_753
timestamp 1644511149
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_765
timestamp 1644511149
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1644511149
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1644511149
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_785
timestamp 1644511149
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_797
timestamp 1644511149
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_809
timestamp 1644511149
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_821
timestamp 1644511149
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1644511149
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1644511149
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_841
timestamp 1644511149
transform 1 0 78476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_495
timestamp 1644511149
transform 1 0 46644 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_500
timestamp 1644511149
transform 1 0 47104 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_524
timestamp 1644511149
transform 1 0 49312 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_713
timestamp 1644511149
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_725
timestamp 1644511149
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_737
timestamp 1644511149
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1644511149
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1644511149
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_757
timestamp 1644511149
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_769
timestamp 1644511149
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_781
timestamp 1644511149
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_793
timestamp 1644511149
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1644511149
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1644511149
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_813
timestamp 1644511149
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_825
timestamp 1644511149
transform 1 0 77004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_829
timestamp 1644511149
transform 1 0 77372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_832
timestamp 1644511149
transform 1 0 77648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_838
timestamp 1644511149
transform 1 0 78200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_525
timestamp 1644511149
transform 1 0 49404 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_530
timestamp 1644511149
transform 1 0 49864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_542
timestamp 1644511149
transform 1 0 50968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_554
timestamp 1644511149
transform 1 0 52072 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1644511149
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_741
timestamp 1644511149
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_753
timestamp 1644511149
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_765
timestamp 1644511149
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1644511149
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1644511149
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_785
timestamp 1644511149
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_797
timestamp 1644511149
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_809
timestamp 1644511149
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_821
timestamp 1644511149
transform 1 0 76636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_827
timestamp 1644511149
transform 1 0 77188 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_830
timestamp 1644511149
transform 1 0 77464 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_836
timestamp 1644511149
transform 1 0 78016 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_841
timestamp 1644511149
transform 1 0 78476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_521
timestamp 1644511149
transform 1 0 49036 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_526
timestamp 1644511149
transform 1 0 49496 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_737
timestamp 1644511149
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1644511149
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1644511149
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_757
timestamp 1644511149
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_769
timestamp 1644511149
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_781
timestamp 1644511149
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_793
timestamp 1644511149
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1644511149
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1644511149
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_813
timestamp 1644511149
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_825
timestamp 1644511149
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_837
timestamp 1644511149
transform 1 0 78108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_841
timestamp 1644511149
transform 1 0 78476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_513
timestamp 1644511149
transform 1 0 48300 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_524
timestamp 1644511149
transform 1 0 49312 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_536
timestamp 1644511149
transform 1 0 50416 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_548
timestamp 1644511149
transform 1 0 51520 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_741
timestamp 1644511149
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_753
timestamp 1644511149
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_765
timestamp 1644511149
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1644511149
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1644511149
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_785
timestamp 1644511149
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_797
timestamp 1644511149
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_809
timestamp 1644511149
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_821
timestamp 1644511149
transform 1 0 76636 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_829
timestamp 1644511149
transform 1 0 77372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_836
timestamp 1644511149
transform 1 0 78016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_841
timestamp 1644511149
transform 1 0 78476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_542
timestamp 1644511149
transform 1 0 50968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_550
timestamp 1644511149
transform 1 0 51704 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_562
timestamp 1644511149
transform 1 0 52808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_574
timestamp 1644511149
transform 1 0 53912 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_586
timestamp 1644511149
transform 1 0 55016 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_737
timestamp 1644511149
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1644511149
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1644511149
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_757
timestamp 1644511149
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_769
timestamp 1644511149
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_781
timestamp 1644511149
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_793
timestamp 1644511149
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1644511149
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1644511149
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_813
timestamp 1644511149
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_825
timestamp 1644511149
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_837
timestamp 1644511149
transform 1 0 78108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_841
timestamp 1644511149
transform 1 0 78476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_629
timestamp 1644511149
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_641
timestamp 1644511149
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_653
timestamp 1644511149
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1644511149
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_741
timestamp 1644511149
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_753
timestamp 1644511149
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_765
timestamp 1644511149
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1644511149
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1644511149
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_785
timestamp 1644511149
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_797
timestamp 1644511149
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_809
timestamp 1644511149
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_821
timestamp 1644511149
transform 1 0 76636 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_829
timestamp 1644511149
transform 1 0 77372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_836
timestamp 1644511149
transform 1 0 78016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_841
timestamp 1644511149
transform 1 0 78476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_553
timestamp 1644511149
transform 1 0 51980 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_563
timestamp 1644511149
transform 1 0 52900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_571
timestamp 1644511149
transform 1 0 53636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_583
timestamp 1644511149
transform 1 0 54740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_625
timestamp 1644511149
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1644511149
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1644511149
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_737
timestamp 1644511149
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1644511149
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1644511149
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_757
timestamp 1644511149
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_769
timestamp 1644511149
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_781
timestamp 1644511149
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_793
timestamp 1644511149
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1644511149
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1644511149
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_813
timestamp 1644511149
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_825
timestamp 1644511149
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_837
timestamp 1644511149
transform 1 0 78108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_841
timestamp 1644511149
transform 1 0 78476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_629
timestamp 1644511149
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_641
timestamp 1644511149
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_653
timestamp 1644511149
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1644511149
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1644511149
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_741
timestamp 1644511149
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_753
timestamp 1644511149
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_765
timestamp 1644511149
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1644511149
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1644511149
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_785
timestamp 1644511149
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_797
timestamp 1644511149
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_809
timestamp 1644511149
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_821
timestamp 1644511149
transform 1 0 76636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_829
timestamp 1644511149
transform 1 0 77372 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_836
timestamp 1644511149
transform 1 0 78016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_841
timestamp 1644511149
transform 1 0 78476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_584
timestamp 1644511149
transform 1 0 54832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_602
timestamp 1644511149
transform 1 0 56488 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_614
timestamp 1644511149
transform 1 0 57592 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_626
timestamp 1644511149
transform 1 0 58696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_638
timestamp 1644511149
transform 1 0 59800 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1644511149
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1644511149
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1644511149
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1644511149
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_737
timestamp 1644511149
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1644511149
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1644511149
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_757
timestamp 1644511149
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_769
timestamp 1644511149
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_781
timestamp 1644511149
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_793
timestamp 1644511149
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1644511149
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1644511149
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_813
timestamp 1644511149
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_825
timestamp 1644511149
transform 1 0 77004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_833
timestamp 1644511149
transform 1 0 77740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_838
timestamp 1644511149
transform 1 0 78200 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_603
timestamp 1644511149
transform 1 0 56580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_653
timestamp 1644511149
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1644511149
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1644511149
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_741
timestamp 1644511149
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_753
timestamp 1644511149
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_765
timestamp 1644511149
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1644511149
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1644511149
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_785
timestamp 1644511149
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_797
timestamp 1644511149
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_809
timestamp 1644511149
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_821
timestamp 1644511149
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_833
timestamp 1644511149
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_839
timestamp 1644511149
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_841
timestamp 1644511149
transform 1 0 78476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1644511149
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1644511149
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1644511149
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1644511149
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1644511149
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_737
timestamp 1644511149
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1644511149
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1644511149
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_757
timestamp 1644511149
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_769
timestamp 1644511149
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_781
timestamp 1644511149
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_793
timestamp 1644511149
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1644511149
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1644511149
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_813
timestamp 1644511149
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_825
timestamp 1644511149
transform 1 0 77004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_833
timestamp 1644511149
transform 1 0 77740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_838
timestamp 1644511149
transform 1 0 78200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_741
timestamp 1644511149
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_753
timestamp 1644511149
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_765
timestamp 1644511149
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1644511149
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1644511149
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_785
timestamp 1644511149
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_797
timestamp 1644511149
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_809
timestamp 1644511149
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_821
timestamp 1644511149
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_833
timestamp 1644511149
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_839
timestamp 1644511149
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_841
timestamp 1644511149
transform 1 0 78476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_636
timestamp 1644511149
transform 1 0 59616 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_654
timestamp 1644511149
transform 1 0 61272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_666
timestamp 1644511149
transform 1 0 62376 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_678
timestamp 1644511149
transform 1 0 63480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_690
timestamp 1644511149
transform 1 0 64584 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_698
timestamp 1644511149
transform 1 0 65320 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_737
timestamp 1644511149
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1644511149
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1644511149
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_757
timestamp 1644511149
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_769
timestamp 1644511149
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_781
timestamp 1644511149
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_793
timestamp 1644511149
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1644511149
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1644511149
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_813
timestamp 1644511149
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_825
timestamp 1644511149
transform 1 0 77004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_833
timestamp 1644511149
transform 1 0 77740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_838
timestamp 1644511149
transform 1 0 78200 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_628
timestamp 1644511149
transform 1 0 58880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_640
timestamp 1644511149
transform 1 0 59984 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_653
timestamp 1644511149
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1644511149
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_741
timestamp 1644511149
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_753
timestamp 1644511149
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_765
timestamp 1644511149
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1644511149
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1644511149
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_785
timestamp 1644511149
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_797
timestamp 1644511149
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_809
timestamp 1644511149
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_821
timestamp 1644511149
transform 1 0 76636 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_829
timestamp 1644511149
transform 1 0 77372 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_836
timestamp 1644511149
transform 1 0 78016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_841
timestamp 1644511149
transform 1 0 78476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1644511149
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_645
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_657
timestamp 1644511149
transform 1 0 61548 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_673
timestamp 1644511149
transform 1 0 63020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_685
timestamp 1644511149
transform 1 0 64124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_697
timestamp 1644511149
transform 1 0 65228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_737
timestamp 1644511149
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1644511149
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1644511149
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_757
timestamp 1644511149
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_769
timestamp 1644511149
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_781
timestamp 1644511149
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_793
timestamp 1644511149
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1644511149
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1644511149
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_813
timestamp 1644511149
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1644511149
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_837
timestamp 1644511149
transform 1 0 78108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_841
timestamp 1644511149
transform 1 0 78476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_666
timestamp 1644511149
transform 1 0 62376 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_677
timestamp 1644511149
transform 1 0 63388 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_687
timestamp 1644511149
transform 1 0 64308 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_699
timestamp 1644511149
transform 1 0 65412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_711
timestamp 1644511149
transform 1 0 66516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_723
timestamp 1644511149
transform 1 0 67620 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1644511149
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_741
timestamp 1644511149
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_753
timestamp 1644511149
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_765
timestamp 1644511149
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1644511149
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1644511149
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_785
timestamp 1644511149
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_797
timestamp 1644511149
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_809
timestamp 1644511149
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_821
timestamp 1644511149
transform 1 0 76636 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_829
timestamp 1644511149
transform 1 0 77372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_836
timestamp 1644511149
transform 1 0 78016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_841
timestamp 1644511149
transform 1 0 78476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_674
timestamp 1644511149
transform 1 0 63112 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_682
timestamp 1644511149
transform 1 0 63848 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_694
timestamp 1644511149
transform 1 0 64952 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_710
timestamp 1644511149
transform 1 0 66424 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_722
timestamp 1644511149
transform 1 0 67528 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_734
timestamp 1644511149
transform 1 0 68632 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_746
timestamp 1644511149
transform 1 0 69736 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_754
timestamp 1644511149
transform 1 0 70472 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_757
timestamp 1644511149
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_769
timestamp 1644511149
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_781
timestamp 1644511149
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_793
timestamp 1644511149
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1644511149
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1644511149
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_813
timestamp 1644511149
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_825
timestamp 1644511149
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_837
timestamp 1644511149
transform 1 0 78108 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_841
timestamp 1644511149
transform 1 0 78476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_706
timestamp 1644511149
transform 1 0 66056 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_718
timestamp 1644511149
transform 1 0 67160 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_726
timestamp 1644511149
transform 1 0 67896 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_741
timestamp 1644511149
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_753
timestamp 1644511149
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_765
timestamp 1644511149
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1644511149
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1644511149
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_785
timestamp 1644511149
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_797
timestamp 1644511149
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_809
timestamp 1644511149
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_821
timestamp 1644511149
transform 1 0 76636 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_829
timestamp 1644511149
transform 1 0 77372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_836
timestamp 1644511149
transform 1 0 78016 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_841
timestamp 1644511149
transform 1 0 78476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_625
timestamp 1644511149
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1644511149
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1644511149
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_713
timestamp 1644511149
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_725
timestamp 1644511149
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_737
timestamp 1644511149
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1644511149
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1644511149
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_757
timestamp 1644511149
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_769
timestamp 1644511149
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_781
timestamp 1644511149
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_793
timestamp 1644511149
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1644511149
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1644511149
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_813
timestamp 1644511149
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_825
timestamp 1644511149
transform 1 0 77004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_833
timestamp 1644511149
transform 1 0 77740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_838
timestamp 1644511149
transform 1 0 78200 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1644511149
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_733
timestamp 1644511149
transform 1 0 68540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_745
timestamp 1644511149
transform 1 0 69644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_757
timestamp 1644511149
transform 1 0 70748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_769
timestamp 1644511149
transform 1 0 71852 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_774
timestamp 1644511149
transform 1 0 72312 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_782
timestamp 1644511149
transform 1 0 73048 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_785
timestamp 1644511149
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_797
timestamp 1644511149
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_809
timestamp 1644511149
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_821
timestamp 1644511149
transform 1 0 76636 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_836
timestamp 1644511149
transform 1 0 78016 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_841
timestamp 1644511149
transform 1 0 78476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_625
timestamp 1644511149
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1644511149
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1644511149
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_721
timestamp 1644511149
transform 1 0 67436 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_733
timestamp 1644511149
transform 1 0 68540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_745
timestamp 1644511149
transform 1 0 69644 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_753
timestamp 1644511149
transform 1 0 70380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_757
timestamp 1644511149
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_769
timestamp 1644511149
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_781
timestamp 1644511149
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_793
timestamp 1644511149
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1644511149
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1644511149
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_813
timestamp 1644511149
transform 1 0 75900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_819
timestamp 1644511149
transform 1 0 76452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_832
timestamp 1644511149
transform 1 0 77648 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_840
timestamp 1644511149
transform 1 0 78384 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1644511149
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1644511149
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_737
timestamp 1644511149
transform 1 0 68908 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_749
timestamp 1644511149
transform 1 0 70012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_756
timestamp 1644511149
transform 1 0 70656 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_768
timestamp 1644511149
transform 1 0 71760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_780
timestamp 1644511149
transform 1 0 72864 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_785
timestamp 1644511149
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_797
timestamp 1644511149
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_809
timestamp 1644511149
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_821
timestamp 1644511149
transform 1 0 76636 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_828
timestamp 1644511149
transform 1 0 77280 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_836
timestamp 1644511149
transform 1 0 78016 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_841
timestamp 1644511149
transform 1 0 78476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_725
timestamp 1644511149
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_737
timestamp 1644511149
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 1644511149
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 1644511149
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_757
timestamp 1644511149
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_769
timestamp 1644511149
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_781
timestamp 1644511149
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_793
timestamp 1644511149
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1644511149
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1644511149
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_813
timestamp 1644511149
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_825
timestamp 1644511149
transform 1 0 77004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_833
timestamp 1644511149
transform 1 0 77740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_838
timestamp 1644511149
transform 1 0 78200 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1644511149
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1644511149
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1644511149
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_741
timestamp 1644511149
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_753
timestamp 1644511149
transform 1 0 70380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_770
timestamp 1644511149
transform 1 0 71944 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 1644511149
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 1644511149
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_785
timestamp 1644511149
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_797
timestamp 1644511149
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_809
timestamp 1644511149
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_821
timestamp 1644511149
transform 1 0 76636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_836
timestamp 1644511149
transform 1 0 78016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_841
timestamp 1644511149
transform 1 0 78476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_713
timestamp 1644511149
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_725
timestamp 1644511149
transform 1 0 67804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_737
timestamp 1644511149
transform 1 0 68908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1644511149
transform 1 0 70012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1644511149
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_757
timestamp 1644511149
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_769
timestamp 1644511149
transform 1 0 71852 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_781
timestamp 1644511149
transform 1 0 72956 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_787
timestamp 1644511149
transform 1 0 73508 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_791
timestamp 1644511149
transform 1 0 73876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_803
timestamp 1644511149
transform 1 0 74980 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1644511149
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_813
timestamp 1644511149
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_825
timestamp 1644511149
transform 1 0 77004 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_830
timestamp 1644511149
transform 1 0 77464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_838
timestamp 1644511149
transform 1 0 78200 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_433
timestamp 1644511149
transform 1 0 40940 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1644511149
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1644511149
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1644511149
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1644511149
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1644511149
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_741
timestamp 1644511149
transform 1 0 69276 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_753
timestamp 1644511149
transform 1 0 70380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_765
timestamp 1644511149
transform 1 0 71484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1644511149
transform 1 0 72588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1644511149
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_794
timestamp 1644511149
transform 1 0 74152 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_809
timestamp 1644511149
transform 1 0 75532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_821
timestamp 1644511149
transform 1 0 76636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_828
timestamp 1644511149
transform 1 0 77280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_836
timestamp 1644511149
transform 1 0 78016 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_841
timestamp 1644511149
transform 1 0 78476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1644511149
transform 1 0 5152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_89
timestamp 1644511149
transform 1 0 9292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_101
timestamp 1644511149
transform 1 0 10396 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_106
timestamp 1644511149
transform 1 0 10856 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_127
timestamp 1644511149
transform 1 0 12788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_148
timestamp 1644511149
transform 1 0 14720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1644511149
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_210
timestamp 1644511149
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1644511149
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_242
timestamp 1644511149
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1644511149
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_257
timestamp 1644511149
transform 1 0 24748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_319
timestamp 1644511149
transform 1 0 30452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_331
timestamp 1644511149
transform 1 0 31556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1644511149
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_347
timestamp 1644511149
transform 1 0 33028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 1644511149
transform 1 0 34132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_381
timestamp 1644511149
transform 1 0 36156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_415
timestamp 1644511149
transform 1 0 39284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_431
timestamp 1644511149
transform 1 0 40756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_443
timestamp 1644511149
transform 1 0 41860 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_447
timestamp 1644511149
transform 1 0 42228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_449
timestamp 1644511149
transform 1 0 42412 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_453
timestamp 1644511149
transform 1 0 42780 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_464
timestamp 1644511149
transform 1 0 43792 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_487
timestamp 1644511149
transform 1 0 45908 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_495
timestamp 1644511149
transform 1 0 46644 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_499
timestamp 1644511149
transform 1 0 47012 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_503
timestamp 1644511149
transform 1 0 47380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_505
timestamp 1644511149
transform 1 0 47564 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_519
timestamp 1644511149
transform 1 0 48852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_540
timestamp 1644511149
transform 1 0 50784 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_552
timestamp 1644511149
transform 1 0 51888 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_564
timestamp 1644511149
transform 1 0 52992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_576
timestamp 1644511149
transform 1 0 54096 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_582
timestamp 1644511149
transform 1 0 54648 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_597
timestamp 1644511149
transform 1 0 56028 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_602
timestamp 1644511149
transform 1 0 56488 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_614
timestamp 1644511149
transform 1 0 57592 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_617
timestamp 1644511149
transform 1 0 57868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_623
timestamp 1644511149
transform 1 0 58420 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_635
timestamp 1644511149
transform 1 0 59524 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1644511149
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_648
timestamp 1644511149
transform 1 0 60720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_660
timestamp 1644511149
transform 1 0 61824 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_664
timestamp 1644511149
transform 1 0 62192 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_673
timestamp 1644511149
transform 1 0 63020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_681
timestamp 1644511149
transform 1 0 63756 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_685
timestamp 1644511149
transform 1 0 64124 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 1644511149
transform 1 0 65228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_706
timestamp 1644511149
transform 1 0 66056 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_718
timestamp 1644511149
transform 1 0 67160 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_726
timestamp 1644511149
transform 1 0 67896 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_732
timestamp 1644511149
transform 1 0 68448 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_747
timestamp 1644511149
transform 1 0 69828 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_755
timestamp 1644511149
transform 1 0 70564 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_757
timestamp 1644511149
transform 1 0 70748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_768
timestamp 1644511149
transform 1 0 71760 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_780
timestamp 1644511149
transform 1 0 72864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_785
timestamp 1644511149
transform 1 0 73324 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_789
timestamp 1644511149
transform 1 0 73692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_801
timestamp 1644511149
transform 1 0 74796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_808
timestamp 1644511149
transform 1 0 75440 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_816
timestamp 1644511149
transform 1 0 76176 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_828
timestamp 1644511149
transform 1 0 77280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_836
timestamp 1644511149
transform 1 0 78016 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_841
timestamp 1644511149
transform 1 0 78476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 78844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 78844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 78844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 78844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 78844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 78844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 78844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 78844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 78844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 78844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 78844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 78844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 78844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 78844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 78844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 78844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 78844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 78844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 78844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 78844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 78844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 78844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 78844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 78844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 78844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 78844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 78844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 78844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 78844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 78844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 78844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 78844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 78844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 78844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 78844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 78844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 78844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 78844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 78844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 78844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 78844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 78844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 78844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 78844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 78844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 78844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 78844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 78844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 78844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 78844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 78844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 78844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 78844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 78844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 78844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 78844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 78844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 78844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 78844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 78844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 78844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 78844 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 78844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 78844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 78844 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 62928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 68080 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 73232 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 78384 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _064_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 49864 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _065_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _066_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _067_
timestamp 1644511149
transform 1 0 23276 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _069_
timestamp 1644511149
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 1644511149
transform 1 0 23092 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _071_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 1644511149
transform 1 0 25392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _073_
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1644511149
transform 1 0 27140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _075_
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _076_
timestamp 1644511149
transform 1 0 36432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _077_
timestamp 1644511149
transform 1 0 29532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _078_
timestamp 1644511149
transform 1 0 30176 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _079_
timestamp 1644511149
transform 1 0 31096 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _080_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _081_
timestamp 1644511149
transform 1 0 33028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _082_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 1644511149
transform 1 0 34868 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1644511149
transform 1 0 36064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _085_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1644511149
transform 1 0 37168 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _087_
timestamp 1644511149
transform 1 0 40112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1644511149
transform 1 0 39652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1644511149
transform 1 0 41032 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1644511149
transform 1 0 41216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 1644511149
transform 1 0 42504 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1644511149
transform 1 0 43700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _094_
timestamp 1644511149
transform 1 0 44436 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 1644511149
transform 1 0 46184 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1644511149
transform 1 0 46736 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1644511149
transform 1 0 49496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1644511149
transform 1 0 48484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _100_
timestamp 1644511149
transform 1 0 49128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1644511149
transform 1 0 51336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 1644511149
transform 1 0 52072 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1644511149
transform 1 0 53268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp 1644511149
transform 1 0 54004 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1644511149
transform 1 0 54556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1644511149
transform 1 0 55660 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1644511149
transform 1 0 56212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1644511149
transform 1 0 62744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1644511149
transform 1 0 58052 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 58696 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1644511149
transform 1 0 60260 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 1644511149
transform 1 0 61548 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _115_
timestamp 1644511149
transform 1 0 62100 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1644511149
transform 1 0 63480 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1644511149
transform 1 0 64032 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _119_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 65780 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1644511149
transform 1 0 71944 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _121_
timestamp 1644511149
transform 1 0 67712 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1644511149
transform 1 0 68264 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _123_
timestamp 1644511149
transform 1 0 69184 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1644511149
transform 1 0 70380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 1644511149
transform 1 0 71116 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1644511149
transform 1 0 72312 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 1644511149
transform 1 0 73324 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1644511149
transform 1 0 73600 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 1644511149
transform 1 0 74704 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1644511149
transform 1 0 75900 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _131_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1644511149
transform 1 0 76820 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1644511149
transform 1 0 77004 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1644511149
transform 1 0 77188 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1644511149
transform 1 0 76176 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _137_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _138_
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _139_
timestamp 1644511149
transform 1 0 8740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1644511149
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _141_
timestamp 1644511149
transform 1 0 8740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp 1644511149
transform 1 0 7912 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _145_
timestamp 1644511149
transform 1 0 9844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _148_
timestamp 1644511149
transform 1 0 14168 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1644511149
transform 1 0 14168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1644511149
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _152_
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1644511149
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _156_
timestamp 1644511149
transform 1 0 14168 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _157_
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _159_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1644511149
transform 1 0 9384 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1644511149
transform -1 0 9384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1644511149
transform 1 0 9752 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1644511149
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _170_
timestamp 1644511149
transform -1 0 14812 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1644511149
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 1644511149
transform -1 0 14720 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _174_
timestamp 1644511149
transform -1 0 17112 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _176_
timestamp 1644511149
transform 1 0 17480 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _178_
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 77464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1644511149
transform 1 0 77464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1644511149
transform 1 0 77648 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 77648 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1644511149
transform 1 0 77464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1644511149
transform 1 0 77464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1644511149
transform 1 0 77464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1644511149
transform 1 0 77648 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1644511149
transform 1 0 77648 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1644511149
transform 1 0 77648 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1644511149
transform 1 0 76544 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1644511149
transform 1 0 41032 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1644511149
transform 1 0 42872 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 46736 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 48576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 50508 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 52716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 54372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 56212 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 21896 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 58144 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 61916 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 63848 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 65780 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 68172 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 69552 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 71484 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 73416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 75164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 77188 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 77740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 33396 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1644511149
transform 1 0 35236 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 41032 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1644511149
transform 1 0 42872 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 48852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1644511149
transform 1 0 50508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 54372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1644511149
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 61916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 63848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 65780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 69552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 71484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1644511149
transform 1 0 73416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1644511149
transform 1 0 75072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 76728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 77648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1644511149
transform 1 0 35236 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 4784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 10488 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 12420 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 14352 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 77832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 77648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 77832 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 77832 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 77832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 77648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 77648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 77648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 77648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 77832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 77832 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 77648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 77832 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 77648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 77648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 77648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 77832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 77648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 77832 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 77832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 77648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 77648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 77648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 76912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 76912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 77648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 77832 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 77832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 77832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 77832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 77648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 77648 0 -1 19584
box -38 -48 406 592
<< labels >>
rlabel metal3 s 79200 1232 80000 1352 6 addr[0]
port 0 nsew signal input
rlabel metal3 s 79200 2184 80000 2304 6 addr[1]
port 1 nsew signal input
rlabel metal3 s 79200 3136 80000 3256 6 addr[2]
port 2 nsew signal input
rlabel metal3 s 79200 4088 80000 4208 6 addr[3]
port 3 nsew signal input
rlabel metal3 s 79200 5040 80000 5160 6 addr[4]
port 4 nsew signal input
rlabel metal3 s 79200 5992 80000 6112 6 addr[5]
port 5 nsew signal input
rlabel metal3 s 79200 6808 80000 6928 6 addr[6]
port 6 nsew signal input
rlabel metal3 s 79200 7760 80000 7880 6 addr[7]
port 7 nsew signal input
rlabel metal3 s 79200 8712 80000 8832 6 addr[8]
port 8 nsew signal input
rlabel metal3 s 79200 9664 80000 9784 6 addr[9]
port 9 nsew signal input
rlabel metal2 s 2778 39200 2834 40000 6 addr_mem0[0]
port 10 nsew signal tristate
rlabel metal2 s 4710 39200 4766 40000 6 addr_mem0[1]
port 11 nsew signal tristate
rlabel metal2 s 6642 39200 6698 40000 6 addr_mem0[2]
port 12 nsew signal tristate
rlabel metal2 s 8482 39200 8538 40000 6 addr_mem0[3]
port 13 nsew signal tristate
rlabel metal2 s 10414 39200 10470 40000 6 addr_mem0[4]
port 14 nsew signal tristate
rlabel metal2 s 12346 39200 12402 40000 6 addr_mem0[5]
port 15 nsew signal tristate
rlabel metal2 s 14278 39200 14334 40000 6 addr_mem0[6]
port 16 nsew signal tristate
rlabel metal2 s 16118 39200 16174 40000 6 addr_mem0[7]
port 17 nsew signal tristate
rlabel metal2 s 18050 39200 18106 40000 6 addr_mem0[8]
port 18 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 addr_mem1[0]
port 19 nsew signal tristate
rlabel metal2 s 4710 0 4766 800 6 addr_mem1[1]
port 20 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 addr_mem1[2]
port 21 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 addr_mem1[3]
port 22 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 addr_mem1[4]
port 23 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 addr_mem1[5]
port 24 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 addr_mem1[6]
port 25 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 addr_mem1[7]
port 26 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 addr_mem1[8]
port 27 nsew signal tristate
rlabel metal3 s 79200 416 80000 536 6 csb
port 28 nsew signal input
rlabel metal2 s 938 39200 994 40000 6 csb_mem0
port 29 nsew signal tristate
rlabel metal2 s 938 0 994 800 6 csb_mem1
port 30 nsew signal tristate
rlabel metal3 s 79200 10616 80000 10736 6 dout[0]
port 31 nsew signal tristate
rlabel metal3 s 79200 19864 80000 19984 6 dout[10]
port 32 nsew signal tristate
rlabel metal3 s 79200 20816 80000 20936 6 dout[11]
port 33 nsew signal tristate
rlabel metal3 s 79200 21768 80000 21888 6 dout[12]
port 34 nsew signal tristate
rlabel metal3 s 79200 22720 80000 22840 6 dout[13]
port 35 nsew signal tristate
rlabel metal3 s 79200 23536 80000 23656 6 dout[14]
port 36 nsew signal tristate
rlabel metal3 s 79200 24488 80000 24608 6 dout[15]
port 37 nsew signal tristate
rlabel metal3 s 79200 25440 80000 25560 6 dout[16]
port 38 nsew signal tristate
rlabel metal3 s 79200 26392 80000 26512 6 dout[17]
port 39 nsew signal tristate
rlabel metal3 s 79200 27344 80000 27464 6 dout[18]
port 40 nsew signal tristate
rlabel metal3 s 79200 28296 80000 28416 6 dout[19]
port 41 nsew signal tristate
rlabel metal3 s 79200 11568 80000 11688 6 dout[1]
port 42 nsew signal tristate
rlabel metal3 s 79200 29112 80000 29232 6 dout[20]
port 43 nsew signal tristate
rlabel metal3 s 79200 30064 80000 30184 6 dout[21]
port 44 nsew signal tristate
rlabel metal3 s 79200 31016 80000 31136 6 dout[22]
port 45 nsew signal tristate
rlabel metal3 s 79200 31968 80000 32088 6 dout[23]
port 46 nsew signal tristate
rlabel metal3 s 79200 32920 80000 33040 6 dout[24]
port 47 nsew signal tristate
rlabel metal3 s 79200 33872 80000 33992 6 dout[25]
port 48 nsew signal tristate
rlabel metal3 s 79200 34688 80000 34808 6 dout[26]
port 49 nsew signal tristate
rlabel metal3 s 79200 35640 80000 35760 6 dout[27]
port 50 nsew signal tristate
rlabel metal3 s 79200 36592 80000 36712 6 dout[28]
port 51 nsew signal tristate
rlabel metal3 s 79200 37544 80000 37664 6 dout[29]
port 52 nsew signal tristate
rlabel metal3 s 79200 12384 80000 12504 6 dout[2]
port 53 nsew signal tristate
rlabel metal3 s 79200 38496 80000 38616 6 dout[30]
port 54 nsew signal tristate
rlabel metal3 s 79200 39448 80000 39568 6 dout[31]
port 55 nsew signal tristate
rlabel metal3 s 79200 13336 80000 13456 6 dout[3]
port 56 nsew signal tristate
rlabel metal3 s 79200 14288 80000 14408 6 dout[4]
port 57 nsew signal tristate
rlabel metal3 s 79200 15240 80000 15360 6 dout[5]
port 58 nsew signal tristate
rlabel metal3 s 79200 16192 80000 16312 6 dout[6]
port 59 nsew signal tristate
rlabel metal3 s 79200 17144 80000 17264 6 dout[7]
port 60 nsew signal tristate
rlabel metal3 s 79200 17960 80000 18080 6 dout[8]
port 61 nsew signal tristate
rlabel metal3 s 79200 18912 80000 19032 6 dout[9]
port 62 nsew signal tristate
rlabel metal2 s 19982 39200 20038 40000 6 dout_mem0[0]
port 63 nsew signal input
rlabel metal2 s 39026 39200 39082 40000 6 dout_mem0[10]
port 64 nsew signal input
rlabel metal2 s 40958 39200 41014 40000 6 dout_mem0[11]
port 65 nsew signal input
rlabel metal2 s 42798 39200 42854 40000 6 dout_mem0[12]
port 66 nsew signal input
rlabel metal2 s 44730 39200 44786 40000 6 dout_mem0[13]
port 67 nsew signal input
rlabel metal2 s 46662 39200 46718 40000 6 dout_mem0[14]
port 68 nsew signal input
rlabel metal2 s 48502 39200 48558 40000 6 dout_mem0[15]
port 69 nsew signal input
rlabel metal2 s 50434 39200 50490 40000 6 dout_mem0[16]
port 70 nsew signal input
rlabel metal2 s 52366 39200 52422 40000 6 dout_mem0[17]
port 71 nsew signal input
rlabel metal2 s 54298 39200 54354 40000 6 dout_mem0[18]
port 72 nsew signal input
rlabel metal2 s 56138 39200 56194 40000 6 dout_mem0[19]
port 73 nsew signal input
rlabel metal2 s 21822 39200 21878 40000 6 dout_mem0[1]
port 74 nsew signal input
rlabel metal2 s 58070 39200 58126 40000 6 dout_mem0[20]
port 75 nsew signal input
rlabel metal2 s 60002 39200 60058 40000 6 dout_mem0[21]
port 76 nsew signal input
rlabel metal2 s 61842 39200 61898 40000 6 dout_mem0[22]
port 77 nsew signal input
rlabel metal2 s 63774 39200 63830 40000 6 dout_mem0[23]
port 78 nsew signal input
rlabel metal2 s 65706 39200 65762 40000 6 dout_mem0[24]
port 79 nsew signal input
rlabel metal2 s 67638 39200 67694 40000 6 dout_mem0[25]
port 80 nsew signal input
rlabel metal2 s 69478 39200 69534 40000 6 dout_mem0[26]
port 81 nsew signal input
rlabel metal2 s 71410 39200 71466 40000 6 dout_mem0[27]
port 82 nsew signal input
rlabel metal2 s 73342 39200 73398 40000 6 dout_mem0[28]
port 83 nsew signal input
rlabel metal2 s 75182 39200 75238 40000 6 dout_mem0[29]
port 84 nsew signal input
rlabel metal2 s 23754 39200 23810 40000 6 dout_mem0[2]
port 85 nsew signal input
rlabel metal2 s 77114 39200 77170 40000 6 dout_mem0[30]
port 86 nsew signal input
rlabel metal2 s 79046 39200 79102 40000 6 dout_mem0[31]
port 87 nsew signal input
rlabel metal2 s 25686 39200 25742 40000 6 dout_mem0[3]
port 88 nsew signal input
rlabel metal2 s 27618 39200 27674 40000 6 dout_mem0[4]
port 89 nsew signal input
rlabel metal2 s 29458 39200 29514 40000 6 dout_mem0[5]
port 90 nsew signal input
rlabel metal2 s 31390 39200 31446 40000 6 dout_mem0[6]
port 91 nsew signal input
rlabel metal2 s 33322 39200 33378 40000 6 dout_mem0[7]
port 92 nsew signal input
rlabel metal2 s 35162 39200 35218 40000 6 dout_mem0[8]
port 93 nsew signal input
rlabel metal2 s 37094 39200 37150 40000 6 dout_mem0[9]
port 94 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 dout_mem1[0]
port 95 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 dout_mem1[10]
port 96 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 dout_mem1[11]
port 97 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 dout_mem1[12]
port 98 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 dout_mem1[13]
port 99 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 dout_mem1[14]
port 100 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 dout_mem1[15]
port 101 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 dout_mem1[16]
port 102 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 dout_mem1[17]
port 103 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 dout_mem1[18]
port 104 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 dout_mem1[19]
port 105 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 dout_mem1[1]
port 106 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 dout_mem1[20]
port 107 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 dout_mem1[21]
port 108 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 dout_mem1[22]
port 109 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 dout_mem1[23]
port 110 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 dout_mem1[24]
port 111 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 dout_mem1[25]
port 112 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 dout_mem1[26]
port 113 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 dout_mem1[27]
port 114 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 dout_mem1[28]
port 115 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 dout_mem1[29]
port 116 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 dout_mem1[2]
port 117 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 dout_mem1[30]
port 118 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 dout_mem1[31]
port 119 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 dout_mem1[3]
port 120 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 dout_mem1[4]
port 121 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 dout_mem1[5]
port 122 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 dout_mem1[6]
port 123 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 dout_mem1[7]
port 124 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 dout_mem1[8]
port 125 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 dout_mem1[9]
port 126 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 128 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 128 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
