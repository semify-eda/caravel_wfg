magic
tech sky130B
magscale 1 2
timestamp 1657806947
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 2128 78844 77840
<< metal2 >>
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17498 0 17554 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19706 0 19762 800
rect 20442 0 20498 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23386 0 23442 800
rect 24122 0 24178 800
rect 24858 0 24914 800
rect 25594 0 25650 800
rect 26330 0 26386 800
rect 27066 0 27122 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 29274 0 29330 800
rect 30010 0 30066 800
rect 30746 0 30802 800
rect 31482 0 31538 800
rect 32218 0 32274 800
rect 32954 0 33010 800
rect 33690 0 33746 800
rect 34426 0 34482 800
rect 35162 0 35218 800
rect 35898 0 35954 800
rect 36634 0 36690 800
rect 37370 0 37426 800
rect 38106 0 38162 800
rect 38842 0 38898 800
rect 39578 0 39634 800
rect 40314 0 40370 800
rect 41050 0 41106 800
rect 41786 0 41842 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 43994 0 44050 800
rect 44730 0 44786 800
rect 45466 0 45522 800
rect 46202 0 46258 800
rect 46938 0 46994 800
rect 47674 0 47730 800
rect 48410 0 48466 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50618 0 50674 800
rect 51354 0 51410 800
rect 52090 0 52146 800
rect 52826 0 52882 800
rect 53562 0 53618 800
rect 54298 0 54354 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59450 0 59506 800
rect 60186 0 60242 800
rect 60922 0 60978 800
rect 61658 0 61714 800
rect 62394 0 62450 800
rect 63130 0 63186 800
rect 63866 0 63922 800
rect 64602 0 64658 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66810 0 66866 800
rect 67546 0 67602 800
rect 68282 0 68338 800
rect 69018 0 69074 800
rect 69754 0 69810 800
rect 70490 0 70546 800
rect 71226 0 71282 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73434 0 73490 800
rect 74170 0 74226 800
rect 74906 0 74962 800
rect 75642 0 75698 800
rect 76378 0 76434 800
rect 77114 0 77170 800
rect 77850 0 77906 800
<< obsm2 >>
rect 1398 856 78182 77829
rect 1398 734 1986 856
rect 2154 734 2722 856
rect 2890 734 3458 856
rect 3626 734 4194 856
rect 4362 734 4930 856
rect 5098 734 5666 856
rect 5834 734 6402 856
rect 6570 734 7138 856
rect 7306 734 7874 856
rect 8042 734 8610 856
rect 8778 734 9346 856
rect 9514 734 10082 856
rect 10250 734 10818 856
rect 10986 734 11554 856
rect 11722 734 12290 856
rect 12458 734 13026 856
rect 13194 734 13762 856
rect 13930 734 14498 856
rect 14666 734 15234 856
rect 15402 734 15970 856
rect 16138 734 16706 856
rect 16874 734 17442 856
rect 17610 734 18178 856
rect 18346 734 18914 856
rect 19082 734 19650 856
rect 19818 734 20386 856
rect 20554 734 21122 856
rect 21290 734 21858 856
rect 22026 734 22594 856
rect 22762 734 23330 856
rect 23498 734 24066 856
rect 24234 734 24802 856
rect 24970 734 25538 856
rect 25706 734 26274 856
rect 26442 734 27010 856
rect 27178 734 27746 856
rect 27914 734 28482 856
rect 28650 734 29218 856
rect 29386 734 29954 856
rect 30122 734 30690 856
rect 30858 734 31426 856
rect 31594 734 32162 856
rect 32330 734 32898 856
rect 33066 734 33634 856
rect 33802 734 34370 856
rect 34538 734 35106 856
rect 35274 734 35842 856
rect 36010 734 36578 856
rect 36746 734 37314 856
rect 37482 734 38050 856
rect 38218 734 38786 856
rect 38954 734 39522 856
rect 39690 734 40258 856
rect 40426 734 40994 856
rect 41162 734 41730 856
rect 41898 734 42466 856
rect 42634 734 43202 856
rect 43370 734 43938 856
rect 44106 734 44674 856
rect 44842 734 45410 856
rect 45578 734 46146 856
rect 46314 734 46882 856
rect 47050 734 47618 856
rect 47786 734 48354 856
rect 48522 734 49090 856
rect 49258 734 49826 856
rect 49994 734 50562 856
rect 50730 734 51298 856
rect 51466 734 52034 856
rect 52202 734 52770 856
rect 52938 734 53506 856
rect 53674 734 54242 856
rect 54410 734 54978 856
rect 55146 734 55714 856
rect 55882 734 56450 856
rect 56618 734 57186 856
rect 57354 734 57922 856
rect 58090 734 58658 856
rect 58826 734 59394 856
rect 59562 734 60130 856
rect 60298 734 60866 856
rect 61034 734 61602 856
rect 61770 734 62338 856
rect 62506 734 63074 856
rect 63242 734 63810 856
rect 63978 734 64546 856
rect 64714 734 65282 856
rect 65450 734 66018 856
rect 66186 734 66754 856
rect 66922 734 67490 856
rect 67658 734 68226 856
rect 68394 734 68962 856
rect 69130 734 69698 856
rect 69866 734 70434 856
rect 70602 734 71170 856
rect 71338 734 71906 856
rect 72074 734 72642 856
rect 72810 734 73378 856
rect 73546 734 74114 856
rect 74282 734 74850 856
rect 75018 734 75586 856
rect 75754 734 76322 856
rect 76490 734 77058 856
rect 77226 734 77794 856
rect 77962 734 78182 856
<< metal3 >>
rect 0 74944 800 75064
rect 79200 74944 80000 75064
rect 0 74264 800 74384
rect 79200 74264 80000 74384
rect 0 73584 800 73704
rect 79200 73584 80000 73704
rect 0 72904 800 73024
rect 79200 72904 80000 73024
rect 0 72224 800 72344
rect 79200 72224 80000 72344
rect 0 71544 800 71664
rect 79200 71544 80000 71664
rect 0 70864 800 70984
rect 79200 70864 80000 70984
rect 0 70184 800 70304
rect 79200 70184 80000 70304
rect 0 69504 800 69624
rect 79200 69504 80000 69624
rect 0 68824 800 68944
rect 79200 68824 80000 68944
rect 0 68144 800 68264
rect 79200 68144 80000 68264
rect 0 67464 800 67584
rect 79200 67464 80000 67584
rect 0 66784 800 66904
rect 79200 66784 80000 66904
rect 0 66104 800 66224
rect 79200 66104 80000 66224
rect 0 65424 800 65544
rect 79200 65424 80000 65544
rect 0 64744 800 64864
rect 79200 64744 80000 64864
rect 0 64064 800 64184
rect 79200 64064 80000 64184
rect 0 63384 800 63504
rect 79200 63384 80000 63504
rect 0 62704 800 62824
rect 79200 62704 80000 62824
rect 0 62024 800 62144
rect 79200 62024 80000 62144
rect 0 61344 800 61464
rect 79200 61344 80000 61464
rect 0 60664 800 60784
rect 79200 60664 80000 60784
rect 0 59984 800 60104
rect 79200 59984 80000 60104
rect 0 59304 800 59424
rect 79200 59304 80000 59424
rect 0 58624 800 58744
rect 79200 58624 80000 58744
rect 0 57944 800 58064
rect 79200 57944 80000 58064
rect 0 57264 800 57384
rect 79200 57264 80000 57384
rect 0 56584 800 56704
rect 79200 56584 80000 56704
rect 0 55904 800 56024
rect 79200 55904 80000 56024
rect 0 55224 800 55344
rect 79200 55224 80000 55344
rect 0 54544 800 54664
rect 79200 54544 80000 54664
rect 0 53864 800 53984
rect 79200 53864 80000 53984
rect 0 53184 800 53304
rect 79200 53184 80000 53304
rect 0 52504 800 52624
rect 79200 52504 80000 52624
rect 0 51824 800 51944
rect 79200 51824 80000 51944
rect 0 51144 800 51264
rect 79200 51144 80000 51264
rect 0 50464 800 50584
rect 79200 50464 80000 50584
rect 0 49784 800 49904
rect 79200 49784 80000 49904
rect 0 49104 800 49224
rect 79200 49104 80000 49224
rect 0 48424 800 48544
rect 79200 48424 80000 48544
rect 0 47744 800 47864
rect 79200 47744 80000 47864
rect 0 47064 800 47184
rect 79200 47064 80000 47184
rect 0 46384 800 46504
rect 79200 46384 80000 46504
rect 0 45704 800 45824
rect 79200 45704 80000 45824
rect 0 45024 800 45144
rect 79200 45024 80000 45144
rect 0 44344 800 44464
rect 79200 44344 80000 44464
rect 0 43664 800 43784
rect 79200 43664 80000 43784
rect 0 42984 800 43104
rect 79200 42984 80000 43104
rect 0 42304 800 42424
rect 79200 42304 80000 42424
rect 0 41624 800 41744
rect 79200 41624 80000 41744
rect 0 40944 800 41064
rect 79200 40944 80000 41064
rect 0 40264 800 40384
rect 79200 40264 80000 40384
rect 0 39584 800 39704
rect 79200 39584 80000 39704
rect 0 38904 800 39024
rect 79200 38904 80000 39024
rect 0 38224 800 38344
rect 79200 38224 80000 38344
rect 0 37544 800 37664
rect 79200 37544 80000 37664
rect 0 36864 800 36984
rect 79200 36864 80000 36984
rect 0 36184 800 36304
rect 79200 36184 80000 36304
rect 0 35504 800 35624
rect 79200 35504 80000 35624
rect 0 34824 800 34944
rect 79200 34824 80000 34944
rect 0 34144 800 34264
rect 79200 34144 80000 34264
rect 0 33464 800 33584
rect 79200 33464 80000 33584
rect 0 32784 800 32904
rect 79200 32784 80000 32904
rect 0 32104 800 32224
rect 79200 32104 80000 32224
rect 0 31424 800 31544
rect 79200 31424 80000 31544
rect 0 30744 800 30864
rect 79200 30744 80000 30864
rect 0 30064 800 30184
rect 79200 30064 80000 30184
rect 0 29384 800 29504
rect 79200 29384 80000 29504
rect 0 28704 800 28824
rect 79200 28704 80000 28824
rect 0 28024 800 28144
rect 79200 28024 80000 28144
rect 0 27344 800 27464
rect 79200 27344 80000 27464
rect 0 26664 800 26784
rect 79200 26664 80000 26784
rect 0 25984 800 26104
rect 79200 25984 80000 26104
rect 0 25304 800 25424
rect 79200 25304 80000 25424
rect 0 24624 800 24744
rect 79200 24624 80000 24744
rect 0 23944 800 24064
rect 79200 23944 80000 24064
rect 0 23264 800 23384
rect 79200 23264 80000 23384
rect 0 22584 800 22704
rect 79200 22584 80000 22704
rect 0 21904 800 22024
rect 79200 21904 80000 22024
rect 0 21224 800 21344
rect 79200 21224 80000 21344
rect 0 20544 800 20664
rect 79200 20544 80000 20664
rect 0 19864 800 19984
rect 79200 19864 80000 19984
rect 0 19184 800 19304
rect 79200 19184 80000 19304
rect 0 18504 800 18624
rect 79200 18504 80000 18624
rect 0 17824 800 17944
rect 79200 17824 80000 17944
rect 0 17144 800 17264
rect 79200 17144 80000 17264
rect 0 16464 800 16584
rect 79200 16464 80000 16584
rect 0 15784 800 15904
rect 79200 15784 80000 15904
rect 0 15104 800 15224
rect 79200 15104 80000 15224
rect 0 14424 800 14544
rect 79200 14424 80000 14544
rect 0 13744 800 13864
rect 79200 13744 80000 13864
rect 0 13064 800 13184
rect 79200 13064 80000 13184
rect 0 12384 800 12504
rect 79200 12384 80000 12504
rect 0 11704 800 11824
rect 79200 11704 80000 11824
rect 0 11024 800 11144
rect 79200 11024 80000 11144
rect 0 10344 800 10464
rect 79200 10344 80000 10464
rect 0 9664 800 9784
rect 79200 9664 80000 9784
rect 0 8984 800 9104
rect 79200 8984 80000 9104
rect 0 8304 800 8424
rect 79200 8304 80000 8424
rect 0 7624 800 7744
rect 79200 7624 80000 7744
rect 0 6944 800 7064
rect 79200 6944 80000 7064
rect 0 6264 800 6384
rect 79200 6264 80000 6384
rect 0 5584 800 5704
rect 79200 5584 80000 5704
rect 0 4904 800 5024
rect 79200 4904 80000 5024
<< obsm3 >>
rect 800 75144 79200 77825
rect 880 74864 79120 75144
rect 800 74464 79200 74864
rect 880 74184 79120 74464
rect 800 73784 79200 74184
rect 880 73504 79120 73784
rect 800 73104 79200 73504
rect 880 72824 79120 73104
rect 800 72424 79200 72824
rect 880 72144 79120 72424
rect 800 71744 79200 72144
rect 880 71464 79120 71744
rect 800 71064 79200 71464
rect 880 70784 79120 71064
rect 800 70384 79200 70784
rect 880 70104 79120 70384
rect 800 69704 79200 70104
rect 880 69424 79120 69704
rect 800 69024 79200 69424
rect 880 68744 79120 69024
rect 800 68344 79200 68744
rect 880 68064 79120 68344
rect 800 67664 79200 68064
rect 880 67384 79120 67664
rect 800 66984 79200 67384
rect 880 66704 79120 66984
rect 800 66304 79200 66704
rect 880 66024 79120 66304
rect 800 65624 79200 66024
rect 880 65344 79120 65624
rect 800 64944 79200 65344
rect 880 64664 79120 64944
rect 800 64264 79200 64664
rect 880 63984 79120 64264
rect 800 63584 79200 63984
rect 880 63304 79120 63584
rect 800 62904 79200 63304
rect 880 62624 79120 62904
rect 800 62224 79200 62624
rect 880 61944 79120 62224
rect 800 61544 79200 61944
rect 880 61264 79120 61544
rect 800 60864 79200 61264
rect 880 60584 79120 60864
rect 800 60184 79200 60584
rect 880 59904 79120 60184
rect 800 59504 79200 59904
rect 880 59224 79120 59504
rect 800 58824 79200 59224
rect 880 58544 79120 58824
rect 800 58144 79200 58544
rect 880 57864 79120 58144
rect 800 57464 79200 57864
rect 880 57184 79120 57464
rect 800 56784 79200 57184
rect 880 56504 79120 56784
rect 800 56104 79200 56504
rect 880 55824 79120 56104
rect 800 55424 79200 55824
rect 880 55144 79120 55424
rect 800 54744 79200 55144
rect 880 54464 79120 54744
rect 800 54064 79200 54464
rect 880 53784 79120 54064
rect 800 53384 79200 53784
rect 880 53104 79120 53384
rect 800 52704 79200 53104
rect 880 52424 79120 52704
rect 800 52024 79200 52424
rect 880 51744 79120 52024
rect 800 51344 79200 51744
rect 880 51064 79120 51344
rect 800 50664 79200 51064
rect 880 50384 79120 50664
rect 800 49984 79200 50384
rect 880 49704 79120 49984
rect 800 49304 79200 49704
rect 880 49024 79120 49304
rect 800 48624 79200 49024
rect 880 48344 79120 48624
rect 800 47944 79200 48344
rect 880 47664 79120 47944
rect 800 47264 79200 47664
rect 880 46984 79120 47264
rect 800 46584 79200 46984
rect 880 46304 79120 46584
rect 800 45904 79200 46304
rect 880 45624 79120 45904
rect 800 45224 79200 45624
rect 880 44944 79120 45224
rect 800 44544 79200 44944
rect 880 44264 79120 44544
rect 800 43864 79200 44264
rect 880 43584 79120 43864
rect 800 43184 79200 43584
rect 880 42904 79120 43184
rect 800 42504 79200 42904
rect 880 42224 79120 42504
rect 800 41824 79200 42224
rect 880 41544 79120 41824
rect 800 41144 79200 41544
rect 880 40864 79120 41144
rect 800 40464 79200 40864
rect 880 40184 79120 40464
rect 800 39784 79200 40184
rect 880 39504 79120 39784
rect 800 39104 79200 39504
rect 880 38824 79120 39104
rect 800 38424 79200 38824
rect 880 38144 79120 38424
rect 800 37744 79200 38144
rect 880 37464 79120 37744
rect 800 37064 79200 37464
rect 880 36784 79120 37064
rect 800 36384 79200 36784
rect 880 36104 79120 36384
rect 800 35704 79200 36104
rect 880 35424 79120 35704
rect 800 35024 79200 35424
rect 880 34744 79120 35024
rect 800 34344 79200 34744
rect 880 34064 79120 34344
rect 800 33664 79200 34064
rect 880 33384 79120 33664
rect 800 32984 79200 33384
rect 880 32704 79120 32984
rect 800 32304 79200 32704
rect 880 32024 79120 32304
rect 800 31624 79200 32024
rect 880 31344 79120 31624
rect 800 30944 79200 31344
rect 880 30664 79120 30944
rect 800 30264 79200 30664
rect 880 29984 79120 30264
rect 800 29584 79200 29984
rect 880 29304 79120 29584
rect 800 28904 79200 29304
rect 880 28624 79120 28904
rect 800 28224 79200 28624
rect 880 27944 79120 28224
rect 800 27544 79200 27944
rect 880 27264 79120 27544
rect 800 26864 79200 27264
rect 880 26584 79120 26864
rect 800 26184 79200 26584
rect 880 25904 79120 26184
rect 800 25504 79200 25904
rect 880 25224 79120 25504
rect 800 24824 79200 25224
rect 880 24544 79120 24824
rect 800 24144 79200 24544
rect 880 23864 79120 24144
rect 800 23464 79200 23864
rect 880 23184 79120 23464
rect 800 22784 79200 23184
rect 880 22504 79120 22784
rect 800 22104 79200 22504
rect 880 21824 79120 22104
rect 800 21424 79200 21824
rect 880 21144 79120 21424
rect 800 20744 79200 21144
rect 880 20464 79120 20744
rect 800 20064 79200 20464
rect 880 19784 79120 20064
rect 800 19384 79200 19784
rect 880 19104 79120 19384
rect 800 18704 79200 19104
rect 880 18424 79120 18704
rect 800 18024 79200 18424
rect 880 17744 79120 18024
rect 800 17344 79200 17744
rect 880 17064 79120 17344
rect 800 16664 79200 17064
rect 880 16384 79120 16664
rect 800 15984 79200 16384
rect 880 15704 79120 15984
rect 800 15304 79200 15704
rect 880 15024 79120 15304
rect 800 14624 79200 15024
rect 880 14344 79120 14624
rect 800 13944 79200 14344
rect 880 13664 79120 13944
rect 800 13264 79200 13664
rect 880 12984 79120 13264
rect 800 12584 79200 12984
rect 880 12304 79120 12584
rect 800 11904 79200 12304
rect 880 11624 79120 11904
rect 800 11224 79200 11624
rect 880 10944 79120 11224
rect 800 10544 79200 10944
rect 880 10264 79120 10544
rect 800 9864 79200 10264
rect 880 9584 79120 9864
rect 800 9184 79200 9584
rect 880 8904 79120 9184
rect 800 8504 79200 8904
rect 880 8224 79120 8504
rect 800 7824 79200 8224
rect 880 7544 79120 7824
rect 800 7144 79200 7544
rect 880 6864 79120 7144
rect 800 6464 79200 6864
rect 880 6184 79120 6464
rect 800 5784 79200 6184
rect 880 5504 79120 5784
rect 800 5104 79200 5504
rect 880 4824 79120 5104
rect 800 2143 79200 4824
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 1715 61099 1781 75309
<< labels >>
rlabel metal2 s 77114 0 77170 800 6 io_wbs_ack
port 1 nsew signal output
rlabel metal3 s 79200 74264 80000 74384 6 io_wbs_ack_0
port 2 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 io_wbs_ack_1
port 3 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 io_wbs_adr[0]
port 4 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 io_wbs_adr[10]
port 5 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 io_wbs_adr[11]
port 6 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_wbs_adr[12]
port 7 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_wbs_adr[13]
port 8 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 io_wbs_adr[14]
port 9 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 io_wbs_adr[15]
port 10 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 io_wbs_adr[16]
port 11 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 io_wbs_adr[17]
port 12 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 io_wbs_adr[18]
port 13 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 io_wbs_adr[19]
port 14 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 io_wbs_adr[1]
port 15 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_adr[20]
port 16 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 io_wbs_adr[21]
port 17 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 io_wbs_adr[22]
port 18 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 io_wbs_adr[23]
port 19 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 io_wbs_adr[24]
port 20 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 io_wbs_adr[25]
port 21 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 io_wbs_adr[26]
port 22 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_wbs_adr[27]
port 23 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 io_wbs_adr[28]
port 24 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 io_wbs_adr[29]
port 25 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 io_wbs_adr[2]
port 26 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 io_wbs_adr[30]
port 27 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 io_wbs_adr[31]
port 28 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 io_wbs_adr[3]
port 29 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 io_wbs_adr[4]
port 30 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 io_wbs_adr[5]
port 31 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_wbs_adr[6]
port 32 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 io_wbs_adr[7]
port 33 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 io_wbs_adr[8]
port 34 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 io_wbs_adr[9]
port 35 nsew signal input
rlabel metal3 s 79200 4904 80000 5024 6 io_wbs_adr_0[0]
port 36 nsew signal output
rlabel metal3 s 79200 11704 80000 11824 6 io_wbs_adr_0[10]
port 37 nsew signal output
rlabel metal3 s 79200 12384 80000 12504 6 io_wbs_adr_0[11]
port 38 nsew signal output
rlabel metal3 s 79200 13064 80000 13184 6 io_wbs_adr_0[12]
port 39 nsew signal output
rlabel metal3 s 79200 13744 80000 13864 6 io_wbs_adr_0[13]
port 40 nsew signal output
rlabel metal3 s 79200 14424 80000 14544 6 io_wbs_adr_0[14]
port 41 nsew signal output
rlabel metal3 s 79200 15104 80000 15224 6 io_wbs_adr_0[15]
port 42 nsew signal output
rlabel metal3 s 79200 15784 80000 15904 6 io_wbs_adr_0[16]
port 43 nsew signal output
rlabel metal3 s 79200 16464 80000 16584 6 io_wbs_adr_0[17]
port 44 nsew signal output
rlabel metal3 s 79200 17144 80000 17264 6 io_wbs_adr_0[18]
port 45 nsew signal output
rlabel metal3 s 79200 17824 80000 17944 6 io_wbs_adr_0[19]
port 46 nsew signal output
rlabel metal3 s 79200 5584 80000 5704 6 io_wbs_adr_0[1]
port 47 nsew signal output
rlabel metal3 s 79200 18504 80000 18624 6 io_wbs_adr_0[20]
port 48 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 io_wbs_adr_0[21]
port 49 nsew signal output
rlabel metal3 s 79200 19864 80000 19984 6 io_wbs_adr_0[22]
port 50 nsew signal output
rlabel metal3 s 79200 20544 80000 20664 6 io_wbs_adr_0[23]
port 51 nsew signal output
rlabel metal3 s 79200 21224 80000 21344 6 io_wbs_adr_0[24]
port 52 nsew signal output
rlabel metal3 s 79200 21904 80000 22024 6 io_wbs_adr_0[25]
port 53 nsew signal output
rlabel metal3 s 79200 22584 80000 22704 6 io_wbs_adr_0[26]
port 54 nsew signal output
rlabel metal3 s 79200 23264 80000 23384 6 io_wbs_adr_0[27]
port 55 nsew signal output
rlabel metal3 s 79200 23944 80000 24064 6 io_wbs_adr_0[28]
port 56 nsew signal output
rlabel metal3 s 79200 24624 80000 24744 6 io_wbs_adr_0[29]
port 57 nsew signal output
rlabel metal3 s 79200 6264 80000 6384 6 io_wbs_adr_0[2]
port 58 nsew signal output
rlabel metal3 s 79200 25304 80000 25424 6 io_wbs_adr_0[30]
port 59 nsew signal output
rlabel metal3 s 79200 25984 80000 26104 6 io_wbs_adr_0[31]
port 60 nsew signal output
rlabel metal3 s 79200 6944 80000 7064 6 io_wbs_adr_0[3]
port 61 nsew signal output
rlabel metal3 s 79200 7624 80000 7744 6 io_wbs_adr_0[4]
port 62 nsew signal output
rlabel metal3 s 79200 8304 80000 8424 6 io_wbs_adr_0[5]
port 63 nsew signal output
rlabel metal3 s 79200 8984 80000 9104 6 io_wbs_adr_0[6]
port 64 nsew signal output
rlabel metal3 s 79200 9664 80000 9784 6 io_wbs_adr_0[7]
port 65 nsew signal output
rlabel metal3 s 79200 10344 80000 10464 6 io_wbs_adr_0[8]
port 66 nsew signal output
rlabel metal3 s 79200 11024 80000 11144 6 io_wbs_adr_0[9]
port 67 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 io_wbs_adr_1[0]
port 68 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 io_wbs_adr_1[10]
port 69 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 io_wbs_adr_1[11]
port 70 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 io_wbs_adr_1[12]
port 71 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 io_wbs_adr_1[13]
port 72 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 io_wbs_adr_1[14]
port 73 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 io_wbs_adr_1[15]
port 74 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 io_wbs_adr_1[16]
port 75 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 io_wbs_adr_1[17]
port 76 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 io_wbs_adr_1[18]
port 77 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 io_wbs_adr_1[19]
port 78 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 io_wbs_adr_1[1]
port 79 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 io_wbs_adr_1[20]
port 80 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 io_wbs_adr_1[21]
port 81 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 io_wbs_adr_1[22]
port 82 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 io_wbs_adr_1[23]
port 83 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 io_wbs_adr_1[24]
port 84 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 io_wbs_adr_1[25]
port 85 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 io_wbs_adr_1[26]
port 86 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 io_wbs_adr_1[27]
port 87 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 io_wbs_adr_1[28]
port 88 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 io_wbs_adr_1[29]
port 89 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 io_wbs_adr_1[2]
port 90 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 io_wbs_adr_1[30]
port 91 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 io_wbs_adr_1[31]
port 92 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 io_wbs_adr_1[3]
port 93 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_wbs_adr_1[4]
port 94 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 io_wbs_adr_1[5]
port 95 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 io_wbs_adr_1[6]
port 96 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 io_wbs_adr_1[7]
port 97 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 io_wbs_adr_1[8]
port 98 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 io_wbs_adr_1[9]
port 99 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 io_wbs_cyc
port 100 nsew signal input
rlabel metal3 s 79200 74944 80000 75064 6 io_wbs_cyc_0
port 101 nsew signal output
rlabel metal3 s 0 74944 800 75064 6 io_wbs_cyc_1
port 102 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 io_wbs_datrd[0]
port 103 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 io_wbs_datrd[10]
port 104 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 io_wbs_datrd[11]
port 105 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 io_wbs_datrd[12]
port 106 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 io_wbs_datrd[13]
port 107 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 io_wbs_datrd[14]
port 108 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 io_wbs_datrd[15]
port 109 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 io_wbs_datrd[16]
port 110 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 io_wbs_datrd[17]
port 111 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 io_wbs_datrd[18]
port 112 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 io_wbs_datrd[19]
port 113 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 io_wbs_datrd[1]
port 114 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 io_wbs_datrd[20]
port 115 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 io_wbs_datrd[21]
port 116 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 io_wbs_datrd[22]
port 117 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 io_wbs_datrd[23]
port 118 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 io_wbs_datrd[24]
port 119 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 io_wbs_datrd[25]
port 120 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 io_wbs_datrd[26]
port 121 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 io_wbs_datrd[27]
port 122 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 io_wbs_datrd[28]
port 123 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 io_wbs_datrd[29]
port 124 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 io_wbs_datrd[2]
port 125 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 io_wbs_datrd[30]
port 126 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 io_wbs_datrd[31]
port 127 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 io_wbs_datrd[3]
port 128 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 io_wbs_datrd[4]
port 129 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 io_wbs_datrd[5]
port 130 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 io_wbs_datrd[6]
port 131 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 io_wbs_datrd[7]
port 132 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 io_wbs_datrd[8]
port 133 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 io_wbs_datrd[9]
port 134 nsew signal output
rlabel metal3 s 79200 48424 80000 48544 6 io_wbs_datrd_0[0]
port 135 nsew signal input
rlabel metal3 s 79200 55224 80000 55344 6 io_wbs_datrd_0[10]
port 136 nsew signal input
rlabel metal3 s 79200 55904 80000 56024 6 io_wbs_datrd_0[11]
port 137 nsew signal input
rlabel metal3 s 79200 56584 80000 56704 6 io_wbs_datrd_0[12]
port 138 nsew signal input
rlabel metal3 s 79200 57264 80000 57384 6 io_wbs_datrd_0[13]
port 139 nsew signal input
rlabel metal3 s 79200 57944 80000 58064 6 io_wbs_datrd_0[14]
port 140 nsew signal input
rlabel metal3 s 79200 58624 80000 58744 6 io_wbs_datrd_0[15]
port 141 nsew signal input
rlabel metal3 s 79200 59304 80000 59424 6 io_wbs_datrd_0[16]
port 142 nsew signal input
rlabel metal3 s 79200 59984 80000 60104 6 io_wbs_datrd_0[17]
port 143 nsew signal input
rlabel metal3 s 79200 60664 80000 60784 6 io_wbs_datrd_0[18]
port 144 nsew signal input
rlabel metal3 s 79200 61344 80000 61464 6 io_wbs_datrd_0[19]
port 145 nsew signal input
rlabel metal3 s 79200 49104 80000 49224 6 io_wbs_datrd_0[1]
port 146 nsew signal input
rlabel metal3 s 79200 62024 80000 62144 6 io_wbs_datrd_0[20]
port 147 nsew signal input
rlabel metal3 s 79200 62704 80000 62824 6 io_wbs_datrd_0[21]
port 148 nsew signal input
rlabel metal3 s 79200 63384 80000 63504 6 io_wbs_datrd_0[22]
port 149 nsew signal input
rlabel metal3 s 79200 64064 80000 64184 6 io_wbs_datrd_0[23]
port 150 nsew signal input
rlabel metal3 s 79200 64744 80000 64864 6 io_wbs_datrd_0[24]
port 151 nsew signal input
rlabel metal3 s 79200 65424 80000 65544 6 io_wbs_datrd_0[25]
port 152 nsew signal input
rlabel metal3 s 79200 66104 80000 66224 6 io_wbs_datrd_0[26]
port 153 nsew signal input
rlabel metal3 s 79200 66784 80000 66904 6 io_wbs_datrd_0[27]
port 154 nsew signal input
rlabel metal3 s 79200 67464 80000 67584 6 io_wbs_datrd_0[28]
port 155 nsew signal input
rlabel metal3 s 79200 68144 80000 68264 6 io_wbs_datrd_0[29]
port 156 nsew signal input
rlabel metal3 s 79200 49784 80000 49904 6 io_wbs_datrd_0[2]
port 157 nsew signal input
rlabel metal3 s 79200 68824 80000 68944 6 io_wbs_datrd_0[30]
port 158 nsew signal input
rlabel metal3 s 79200 69504 80000 69624 6 io_wbs_datrd_0[31]
port 159 nsew signal input
rlabel metal3 s 79200 50464 80000 50584 6 io_wbs_datrd_0[3]
port 160 nsew signal input
rlabel metal3 s 79200 51144 80000 51264 6 io_wbs_datrd_0[4]
port 161 nsew signal input
rlabel metal3 s 79200 51824 80000 51944 6 io_wbs_datrd_0[5]
port 162 nsew signal input
rlabel metal3 s 79200 52504 80000 52624 6 io_wbs_datrd_0[6]
port 163 nsew signal input
rlabel metal3 s 79200 53184 80000 53304 6 io_wbs_datrd_0[7]
port 164 nsew signal input
rlabel metal3 s 79200 53864 80000 53984 6 io_wbs_datrd_0[8]
port 165 nsew signal input
rlabel metal3 s 79200 54544 80000 54664 6 io_wbs_datrd_0[9]
port 166 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 io_wbs_datrd_1[0]
port 167 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 io_wbs_datrd_1[10]
port 168 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 io_wbs_datrd_1[11]
port 169 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 io_wbs_datrd_1[12]
port 170 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 io_wbs_datrd_1[13]
port 171 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 io_wbs_datrd_1[14]
port 172 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 io_wbs_datrd_1[15]
port 173 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 io_wbs_datrd_1[16]
port 174 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 io_wbs_datrd_1[17]
port 175 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 io_wbs_datrd_1[18]
port 176 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 io_wbs_datrd_1[19]
port 177 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 io_wbs_datrd_1[1]
port 178 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 io_wbs_datrd_1[20]
port 179 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 io_wbs_datrd_1[21]
port 180 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 io_wbs_datrd_1[22]
port 181 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 io_wbs_datrd_1[23]
port 182 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_wbs_datrd_1[24]
port 183 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 io_wbs_datrd_1[25]
port 184 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 io_wbs_datrd_1[26]
port 185 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 io_wbs_datrd_1[27]
port 186 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 io_wbs_datrd_1[28]
port 187 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 io_wbs_datrd_1[29]
port 188 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 io_wbs_datrd_1[2]
port 189 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 io_wbs_datrd_1[30]
port 190 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 io_wbs_datrd_1[31]
port 191 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 io_wbs_datrd_1[3]
port 192 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 io_wbs_datrd_1[4]
port 193 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 io_wbs_datrd_1[5]
port 194 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 io_wbs_datrd_1[6]
port 195 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 io_wbs_datrd_1[7]
port 196 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 io_wbs_datrd_1[8]
port 197 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 io_wbs_datrd_1[9]
port 198 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 io_wbs_datwr[0]
port 199 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 io_wbs_datwr[10]
port 200 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 io_wbs_datwr[11]
port 201 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 io_wbs_datwr[12]
port 202 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 io_wbs_datwr[13]
port 203 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 io_wbs_datwr[14]
port 204 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 io_wbs_datwr[15]
port 205 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 io_wbs_datwr[16]
port 206 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 io_wbs_datwr[17]
port 207 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 io_wbs_datwr[18]
port 208 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 io_wbs_datwr[19]
port 209 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 io_wbs_datwr[1]
port 210 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 io_wbs_datwr[20]
port 211 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 io_wbs_datwr[21]
port 212 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 io_wbs_datwr[22]
port 213 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 io_wbs_datwr[23]
port 214 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 io_wbs_datwr[24]
port 215 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 io_wbs_datwr[25]
port 216 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 io_wbs_datwr[26]
port 217 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 io_wbs_datwr[27]
port 218 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 io_wbs_datwr[28]
port 219 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 io_wbs_datwr[29]
port 220 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 io_wbs_datwr[2]
port 221 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_wbs_datwr[30]
port 222 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 io_wbs_datwr[31]
port 223 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 io_wbs_datwr[3]
port 224 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 io_wbs_datwr[4]
port 225 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 io_wbs_datwr[5]
port 226 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 io_wbs_datwr[6]
port 227 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 io_wbs_datwr[7]
port 228 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 io_wbs_datwr[8]
port 229 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 io_wbs_datwr[9]
port 230 nsew signal input
rlabel metal3 s 79200 26664 80000 26784 6 io_wbs_datwr_0[0]
port 231 nsew signal output
rlabel metal3 s 79200 33464 80000 33584 6 io_wbs_datwr_0[10]
port 232 nsew signal output
rlabel metal3 s 79200 34144 80000 34264 6 io_wbs_datwr_0[11]
port 233 nsew signal output
rlabel metal3 s 79200 34824 80000 34944 6 io_wbs_datwr_0[12]
port 234 nsew signal output
rlabel metal3 s 79200 35504 80000 35624 6 io_wbs_datwr_0[13]
port 235 nsew signal output
rlabel metal3 s 79200 36184 80000 36304 6 io_wbs_datwr_0[14]
port 236 nsew signal output
rlabel metal3 s 79200 36864 80000 36984 6 io_wbs_datwr_0[15]
port 237 nsew signal output
rlabel metal3 s 79200 37544 80000 37664 6 io_wbs_datwr_0[16]
port 238 nsew signal output
rlabel metal3 s 79200 38224 80000 38344 6 io_wbs_datwr_0[17]
port 239 nsew signal output
rlabel metal3 s 79200 38904 80000 39024 6 io_wbs_datwr_0[18]
port 240 nsew signal output
rlabel metal3 s 79200 39584 80000 39704 6 io_wbs_datwr_0[19]
port 241 nsew signal output
rlabel metal3 s 79200 27344 80000 27464 6 io_wbs_datwr_0[1]
port 242 nsew signal output
rlabel metal3 s 79200 40264 80000 40384 6 io_wbs_datwr_0[20]
port 243 nsew signal output
rlabel metal3 s 79200 40944 80000 41064 6 io_wbs_datwr_0[21]
port 244 nsew signal output
rlabel metal3 s 79200 41624 80000 41744 6 io_wbs_datwr_0[22]
port 245 nsew signal output
rlabel metal3 s 79200 42304 80000 42424 6 io_wbs_datwr_0[23]
port 246 nsew signal output
rlabel metal3 s 79200 42984 80000 43104 6 io_wbs_datwr_0[24]
port 247 nsew signal output
rlabel metal3 s 79200 43664 80000 43784 6 io_wbs_datwr_0[25]
port 248 nsew signal output
rlabel metal3 s 79200 44344 80000 44464 6 io_wbs_datwr_0[26]
port 249 nsew signal output
rlabel metal3 s 79200 45024 80000 45144 6 io_wbs_datwr_0[27]
port 250 nsew signal output
rlabel metal3 s 79200 45704 80000 45824 6 io_wbs_datwr_0[28]
port 251 nsew signal output
rlabel metal3 s 79200 46384 80000 46504 6 io_wbs_datwr_0[29]
port 252 nsew signal output
rlabel metal3 s 79200 28024 80000 28144 6 io_wbs_datwr_0[2]
port 253 nsew signal output
rlabel metal3 s 79200 47064 80000 47184 6 io_wbs_datwr_0[30]
port 254 nsew signal output
rlabel metal3 s 79200 47744 80000 47864 6 io_wbs_datwr_0[31]
port 255 nsew signal output
rlabel metal3 s 79200 28704 80000 28824 6 io_wbs_datwr_0[3]
port 256 nsew signal output
rlabel metal3 s 79200 29384 80000 29504 6 io_wbs_datwr_0[4]
port 257 nsew signal output
rlabel metal3 s 79200 30064 80000 30184 6 io_wbs_datwr_0[5]
port 258 nsew signal output
rlabel metal3 s 79200 30744 80000 30864 6 io_wbs_datwr_0[6]
port 259 nsew signal output
rlabel metal3 s 79200 31424 80000 31544 6 io_wbs_datwr_0[7]
port 260 nsew signal output
rlabel metal3 s 79200 32104 80000 32224 6 io_wbs_datwr_0[8]
port 261 nsew signal output
rlabel metal3 s 79200 32784 80000 32904 6 io_wbs_datwr_0[9]
port 262 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_wbs_datwr_1[0]
port 263 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 io_wbs_datwr_1[10]
port 264 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 io_wbs_datwr_1[11]
port 265 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 io_wbs_datwr_1[12]
port 266 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 io_wbs_datwr_1[13]
port 267 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 io_wbs_datwr_1[14]
port 268 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 io_wbs_datwr_1[15]
port 269 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 io_wbs_datwr_1[16]
port 270 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 io_wbs_datwr_1[17]
port 271 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 io_wbs_datwr_1[18]
port 272 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 io_wbs_datwr_1[19]
port 273 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 io_wbs_datwr_1[1]
port 274 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 io_wbs_datwr_1[20]
port 275 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_wbs_datwr_1[21]
port 276 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 io_wbs_datwr_1[22]
port 277 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 io_wbs_datwr_1[23]
port 278 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 io_wbs_datwr_1[24]
port 279 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 io_wbs_datwr_1[25]
port 280 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 io_wbs_datwr_1[26]
port 281 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 io_wbs_datwr_1[27]
port 282 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 io_wbs_datwr_1[28]
port 283 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 io_wbs_datwr_1[29]
port 284 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 io_wbs_datwr_1[2]
port 285 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_wbs_datwr_1[30]
port 286 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 io_wbs_datwr_1[31]
port 287 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 io_wbs_datwr_1[3]
port 288 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_wbs_datwr_1[4]
port 289 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 io_wbs_datwr_1[5]
port 290 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 io_wbs_datwr_1[6]
port 291 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 io_wbs_datwr_1[7]
port 292 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 io_wbs_datwr_1[8]
port 293 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 io_wbs_datwr_1[9]
port 294 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 io_wbs_sel[0]
port 295 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 io_wbs_sel[1]
port 296 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 io_wbs_sel[2]
port 297 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 io_wbs_sel[3]
port 298 nsew signal input
rlabel metal3 s 79200 70864 80000 70984 6 io_wbs_sel_0[0]
port 299 nsew signal output
rlabel metal3 s 79200 71544 80000 71664 6 io_wbs_sel_0[1]
port 300 nsew signal output
rlabel metal3 s 79200 72224 80000 72344 6 io_wbs_sel_0[2]
port 301 nsew signal output
rlabel metal3 s 79200 72904 80000 73024 6 io_wbs_sel_0[3]
port 302 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 io_wbs_sel_1[0]
port 303 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 io_wbs_sel_1[1]
port 304 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 io_wbs_sel_1[2]
port 305 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 io_wbs_sel_1[3]
port 306 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 io_wbs_stb
port 307 nsew signal input
rlabel metal3 s 79200 73584 80000 73704 6 io_wbs_stb_0
port 308 nsew signal output
rlabel metal3 s 0 73584 800 73704 6 io_wbs_stb_1
port 309 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 io_wbs_we
port 310 nsew signal input
rlabel metal3 s 79200 70184 80000 70304 6 io_wbs_we_0
port 311 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 io_wbs_we_1
port 312 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 313 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 313 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 313 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 314 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 314 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2751964
string GDS_FILE /home/leo/Dokumente/caravel_workspace_mpw7/caravel_wfg/openlane/wb_mux/runs/22_07_14_15_55/results/signoff/wb_mux.magic.gds
string GDS_START 97368
<< end >>

