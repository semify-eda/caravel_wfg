magic
tech sky130A
magscale 1 2
timestamp 1657176828
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 382 1708 79658 77840
<< metal2 >>
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4342 0 4398 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8390 0 8446 800
rect 9126 0 9182 800
rect 9954 0 10010 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 13910 0 13966 800
rect 14738 0 14794 800
rect 15566 0 15622 800
rect 16394 0 16450 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19522 0 19578 800
rect 20350 0 20406 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22742 0 22798 800
rect 23570 0 23626 800
rect 24398 0 24454 800
rect 25134 0 25190 800
rect 25962 0 26018 800
rect 26790 0 26846 800
rect 27526 0 27582 800
rect 28354 0 28410 800
rect 29182 0 29238 800
rect 29918 0 29974 800
rect 30746 0 30802 800
rect 31574 0 31630 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33966 0 34022 800
rect 34794 0 34850 800
rect 35530 0 35586 800
rect 36358 0 36414 800
rect 37186 0 37242 800
rect 37922 0 37978 800
rect 38750 0 38806 800
rect 39578 0 39634 800
rect 40406 0 40462 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45190 0 45246 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47582 0 47638 800
rect 48410 0 48466 800
rect 49146 0 49202 800
rect 49974 0 50030 800
rect 50802 0 50858 800
rect 51538 0 51594 800
rect 52366 0 52422 800
rect 53194 0 53250 800
rect 53930 0 53986 800
rect 54758 0 54814 800
rect 55586 0 55642 800
rect 56414 0 56470 800
rect 57150 0 57206 800
rect 57978 0 58034 800
rect 58806 0 58862 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61198 0 61254 800
rect 61934 0 61990 800
rect 62762 0 62818 800
rect 63590 0 63646 800
rect 64418 0 64474 800
rect 65154 0 65210 800
rect 65982 0 66038 800
rect 66810 0 66866 800
rect 67546 0 67602 800
rect 68374 0 68430 800
rect 69202 0 69258 800
rect 69938 0 69994 800
rect 70766 0 70822 800
rect 71594 0 71650 800
rect 72422 0 72478 800
rect 73158 0 73214 800
rect 73986 0 74042 800
rect 74814 0 74870 800
rect 75550 0 75606 800
rect 76378 0 76434 800
rect 77206 0 77262 800
rect 77942 0 77998 800
rect 78770 0 78826 800
rect 79598 0 79654 800
<< obsm2 >>
rect 388 856 79652 79529
rect 498 303 1066 856
rect 1234 303 1894 856
rect 2062 303 2722 856
rect 2890 303 3458 856
rect 3626 303 4286 856
rect 4454 303 5114 856
rect 5282 303 5850 856
rect 6018 303 6678 856
rect 6846 303 7506 856
rect 7674 303 8334 856
rect 8502 303 9070 856
rect 9238 303 9898 856
rect 10066 303 10726 856
rect 10894 303 11462 856
rect 11630 303 12290 856
rect 12458 303 13118 856
rect 13286 303 13854 856
rect 14022 303 14682 856
rect 14850 303 15510 856
rect 15678 303 16338 856
rect 16506 303 17074 856
rect 17242 303 17902 856
rect 18070 303 18730 856
rect 18898 303 19466 856
rect 19634 303 20294 856
rect 20462 303 21122 856
rect 21290 303 21858 856
rect 22026 303 22686 856
rect 22854 303 23514 856
rect 23682 303 24342 856
rect 24510 303 25078 856
rect 25246 303 25906 856
rect 26074 303 26734 856
rect 26902 303 27470 856
rect 27638 303 28298 856
rect 28466 303 29126 856
rect 29294 303 29862 856
rect 30030 303 30690 856
rect 30858 303 31518 856
rect 31686 303 32346 856
rect 32514 303 33082 856
rect 33250 303 33910 856
rect 34078 303 34738 856
rect 34906 303 35474 856
rect 35642 303 36302 856
rect 36470 303 37130 856
rect 37298 303 37866 856
rect 38034 303 38694 856
rect 38862 303 39522 856
rect 39690 303 40350 856
rect 40518 303 41086 856
rect 41254 303 41914 856
rect 42082 303 42742 856
rect 42910 303 43478 856
rect 43646 303 44306 856
rect 44474 303 45134 856
rect 45302 303 45870 856
rect 46038 303 46698 856
rect 46866 303 47526 856
rect 47694 303 48354 856
rect 48522 303 49090 856
rect 49258 303 49918 856
rect 50086 303 50746 856
rect 50914 303 51482 856
rect 51650 303 52310 856
rect 52478 303 53138 856
rect 53306 303 53874 856
rect 54042 303 54702 856
rect 54870 303 55530 856
rect 55698 303 56358 856
rect 56526 303 57094 856
rect 57262 303 57922 856
rect 58090 303 58750 856
rect 58918 303 59486 856
rect 59654 303 60314 856
rect 60482 303 61142 856
rect 61310 303 61878 856
rect 62046 303 62706 856
rect 62874 303 63534 856
rect 63702 303 64362 856
rect 64530 303 65098 856
rect 65266 303 65926 856
rect 66094 303 66754 856
rect 66922 303 67490 856
rect 67658 303 68318 856
rect 68486 303 69146 856
rect 69314 303 69882 856
rect 70050 303 70710 856
rect 70878 303 71538 856
rect 71706 303 72366 856
rect 72534 303 73102 856
rect 73270 303 73930 856
rect 74098 303 74758 856
rect 74926 303 75494 856
rect 75662 303 76322 856
rect 76490 303 77150 856
rect 77318 303 77886 856
rect 78054 303 78714 856
rect 78882 303 79542 856
<< metal3 >>
rect 0 79432 800 79552
rect 79200 79432 80000 79552
rect 0 78616 800 78736
rect 79200 78616 80000 78736
rect 0 77800 800 77920
rect 79200 77800 80000 77920
rect 0 76984 800 77104
rect 79200 76984 80000 77104
rect 0 76168 800 76288
rect 79200 76168 80000 76288
rect 0 75352 800 75472
rect 79200 75352 80000 75472
rect 0 74536 800 74656
rect 79200 74536 80000 74656
rect 0 73720 800 73840
rect 79200 73720 80000 73840
rect 0 73040 800 73160
rect 79200 73040 80000 73160
rect 0 72224 800 72344
rect 79200 72224 80000 72344
rect 0 71408 800 71528
rect 79200 71408 80000 71528
rect 0 70592 800 70712
rect 79200 70592 80000 70712
rect 0 69776 800 69896
rect 79200 69776 80000 69896
rect 0 68960 800 69080
rect 79200 68960 80000 69080
rect 0 68144 800 68264
rect 79200 68144 80000 68264
rect 0 67328 800 67448
rect 79200 67328 80000 67448
rect 0 66648 800 66768
rect 79200 66648 80000 66768
rect 0 65832 800 65952
rect 79200 65832 80000 65952
rect 0 65016 800 65136
rect 79200 65016 80000 65136
rect 0 64200 800 64320
rect 79200 64200 80000 64320
rect 0 63384 800 63504
rect 79200 63384 80000 63504
rect 0 62568 800 62688
rect 79200 62568 80000 62688
rect 0 61752 800 61872
rect 79200 61752 80000 61872
rect 0 60936 800 61056
rect 79200 60936 80000 61056
rect 0 60256 800 60376
rect 79200 60256 80000 60376
rect 0 59440 800 59560
rect 79200 59440 80000 59560
rect 0 58624 800 58744
rect 79200 58624 80000 58744
rect 0 57808 800 57928
rect 79200 57808 80000 57928
rect 0 56992 800 57112
rect 79200 56992 80000 57112
rect 0 56176 800 56296
rect 79200 56176 80000 56296
rect 0 55360 800 55480
rect 79200 55360 80000 55480
rect 0 54544 800 54664
rect 79200 54544 80000 54664
rect 0 53728 800 53848
rect 79200 53728 80000 53848
rect 0 53048 800 53168
rect 79200 53048 80000 53168
rect 0 52232 800 52352
rect 79200 52232 80000 52352
rect 0 51416 800 51536
rect 79200 51416 80000 51536
rect 0 50600 800 50720
rect 79200 50600 80000 50720
rect 0 49784 800 49904
rect 79200 49784 80000 49904
rect 0 48968 800 49088
rect 79200 48968 80000 49088
rect 0 48152 800 48272
rect 79200 48152 80000 48272
rect 0 47336 800 47456
rect 79200 47336 80000 47456
rect 0 46656 800 46776
rect 79200 46656 80000 46776
rect 0 45840 800 45960
rect 79200 45840 80000 45960
rect 0 45024 800 45144
rect 79200 45024 80000 45144
rect 0 44208 800 44328
rect 79200 44208 80000 44328
rect 0 43392 800 43512
rect 79200 43392 80000 43512
rect 0 42576 800 42696
rect 79200 42576 80000 42696
rect 0 41760 800 41880
rect 79200 41760 80000 41880
rect 0 40944 800 41064
rect 79200 40944 80000 41064
rect 0 40264 800 40384
rect 79200 40264 80000 40384
rect 0 39448 800 39568
rect 79200 39448 80000 39568
rect 0 38632 800 38752
rect 79200 38632 80000 38752
rect 0 37816 800 37936
rect 79200 37816 80000 37936
rect 0 37000 800 37120
rect 79200 37000 80000 37120
rect 0 36184 800 36304
rect 79200 36184 80000 36304
rect 0 35368 800 35488
rect 79200 35368 80000 35488
rect 0 34552 800 34672
rect 79200 34552 80000 34672
rect 0 33736 800 33856
rect 79200 33736 80000 33856
rect 0 33056 800 33176
rect 79200 33056 80000 33176
rect 0 32240 800 32360
rect 79200 32240 80000 32360
rect 0 31424 800 31544
rect 79200 31424 80000 31544
rect 0 30608 800 30728
rect 79200 30608 80000 30728
rect 0 29792 800 29912
rect 79200 29792 80000 29912
rect 0 28976 800 29096
rect 79200 28976 80000 29096
rect 0 28160 800 28280
rect 79200 28160 80000 28280
rect 0 27344 800 27464
rect 79200 27344 80000 27464
rect 0 26664 800 26784
rect 79200 26664 80000 26784
rect 0 25848 800 25968
rect 79200 25848 80000 25968
rect 0 25032 800 25152
rect 79200 25032 80000 25152
rect 0 24216 800 24336
rect 79200 24216 80000 24336
rect 0 23400 800 23520
rect 79200 23400 80000 23520
rect 0 22584 800 22704
rect 79200 22584 80000 22704
rect 0 21768 800 21888
rect 79200 21768 80000 21888
rect 0 20952 800 21072
rect 79200 20952 80000 21072
rect 0 20272 800 20392
rect 79200 20272 80000 20392
rect 0 19456 800 19576
rect 79200 19456 80000 19576
rect 0 18640 800 18760
rect 79200 18640 80000 18760
rect 0 17824 800 17944
rect 79200 17824 80000 17944
rect 0 17008 800 17128
rect 79200 17008 80000 17128
rect 0 16192 800 16312
rect 79200 16192 80000 16312
rect 0 15376 800 15496
rect 79200 15376 80000 15496
rect 0 14560 800 14680
rect 79200 14560 80000 14680
rect 0 13744 800 13864
rect 79200 13744 80000 13864
rect 0 13064 800 13184
rect 79200 13064 80000 13184
rect 0 12248 800 12368
rect 79200 12248 80000 12368
rect 0 11432 800 11552
rect 79200 11432 80000 11552
rect 0 10616 800 10736
rect 79200 10616 80000 10736
rect 0 9800 800 9920
rect 79200 9800 80000 9920
rect 0 8984 800 9104
rect 79200 8984 80000 9104
rect 0 8168 800 8288
rect 79200 8168 80000 8288
rect 0 7352 800 7472
rect 79200 7352 80000 7472
rect 0 6672 800 6792
rect 79200 6672 80000 6792
rect 0 5856 800 5976
rect 79200 5856 80000 5976
rect 0 5040 800 5160
rect 79200 5040 80000 5160
rect 0 4224 800 4344
rect 79200 4224 80000 4344
rect 0 3408 800 3528
rect 79200 3408 80000 3528
rect 0 2592 800 2712
rect 79200 2592 80000 2712
rect 0 1776 800 1896
rect 79200 1776 80000 1896
rect 0 960 800 1080
rect 79200 960 80000 1080
rect 0 280 800 400
rect 79200 280 80000 400
<< obsm3 >>
rect 880 79352 79120 79525
rect 800 78816 79200 79352
rect 880 78536 79120 78816
rect 800 78000 79200 78536
rect 880 77720 79120 78000
rect 800 77184 79200 77720
rect 880 76904 79120 77184
rect 800 76368 79200 76904
rect 880 76088 79120 76368
rect 800 75552 79200 76088
rect 880 75272 79120 75552
rect 800 74736 79200 75272
rect 880 74456 79120 74736
rect 800 73920 79200 74456
rect 880 73640 79120 73920
rect 800 73240 79200 73640
rect 880 72960 79120 73240
rect 800 72424 79200 72960
rect 880 72144 79120 72424
rect 800 71608 79200 72144
rect 880 71328 79120 71608
rect 800 70792 79200 71328
rect 880 70512 79120 70792
rect 800 69976 79200 70512
rect 880 69696 79120 69976
rect 800 69160 79200 69696
rect 880 68880 79120 69160
rect 800 68344 79200 68880
rect 880 68064 79120 68344
rect 800 67528 79200 68064
rect 880 67248 79120 67528
rect 800 66848 79200 67248
rect 880 66568 79120 66848
rect 800 66032 79200 66568
rect 880 65752 79120 66032
rect 800 65216 79200 65752
rect 880 64936 79120 65216
rect 800 64400 79200 64936
rect 880 64120 79120 64400
rect 800 63584 79200 64120
rect 880 63304 79120 63584
rect 800 62768 79200 63304
rect 880 62488 79120 62768
rect 800 61952 79200 62488
rect 880 61672 79120 61952
rect 800 61136 79200 61672
rect 880 60856 79120 61136
rect 800 60456 79200 60856
rect 880 60176 79120 60456
rect 800 59640 79200 60176
rect 880 59360 79120 59640
rect 800 58824 79200 59360
rect 880 58544 79120 58824
rect 800 58008 79200 58544
rect 880 57728 79120 58008
rect 800 57192 79200 57728
rect 880 56912 79120 57192
rect 800 56376 79200 56912
rect 880 56096 79120 56376
rect 800 55560 79200 56096
rect 880 55280 79120 55560
rect 800 54744 79200 55280
rect 880 54464 79120 54744
rect 800 53928 79200 54464
rect 880 53648 79120 53928
rect 800 53248 79200 53648
rect 880 52968 79120 53248
rect 800 52432 79200 52968
rect 880 52152 79120 52432
rect 800 51616 79200 52152
rect 880 51336 79120 51616
rect 800 50800 79200 51336
rect 880 50520 79120 50800
rect 800 49984 79200 50520
rect 880 49704 79120 49984
rect 800 49168 79200 49704
rect 880 48888 79120 49168
rect 800 48352 79200 48888
rect 880 48072 79120 48352
rect 800 47536 79200 48072
rect 880 47256 79120 47536
rect 800 46856 79200 47256
rect 880 46576 79120 46856
rect 800 46040 79200 46576
rect 880 45760 79120 46040
rect 800 45224 79200 45760
rect 880 44944 79120 45224
rect 800 44408 79200 44944
rect 880 44128 79120 44408
rect 800 43592 79200 44128
rect 880 43312 79120 43592
rect 800 42776 79200 43312
rect 880 42496 79120 42776
rect 800 41960 79200 42496
rect 880 41680 79120 41960
rect 800 41144 79200 41680
rect 880 40864 79120 41144
rect 800 40464 79200 40864
rect 880 40184 79120 40464
rect 800 39648 79200 40184
rect 880 39368 79120 39648
rect 800 38832 79200 39368
rect 880 38552 79120 38832
rect 800 38016 79200 38552
rect 880 37736 79120 38016
rect 800 37200 79200 37736
rect 880 36920 79120 37200
rect 800 36384 79200 36920
rect 880 36104 79120 36384
rect 800 35568 79200 36104
rect 880 35288 79120 35568
rect 800 34752 79200 35288
rect 880 34472 79120 34752
rect 800 33936 79200 34472
rect 880 33656 79120 33936
rect 800 33256 79200 33656
rect 880 32976 79120 33256
rect 800 32440 79200 32976
rect 880 32160 79120 32440
rect 800 31624 79200 32160
rect 880 31344 79120 31624
rect 800 30808 79200 31344
rect 880 30528 79120 30808
rect 800 29992 79200 30528
rect 880 29712 79120 29992
rect 800 29176 79200 29712
rect 880 28896 79120 29176
rect 800 28360 79200 28896
rect 880 28080 79120 28360
rect 800 27544 79200 28080
rect 880 27264 79120 27544
rect 800 26864 79200 27264
rect 880 26584 79120 26864
rect 800 26048 79200 26584
rect 880 25768 79120 26048
rect 800 25232 79200 25768
rect 880 24952 79120 25232
rect 800 24416 79200 24952
rect 880 24136 79120 24416
rect 800 23600 79200 24136
rect 880 23320 79120 23600
rect 800 22784 79200 23320
rect 880 22504 79120 22784
rect 800 21968 79200 22504
rect 880 21688 79120 21968
rect 800 21152 79200 21688
rect 880 20872 79120 21152
rect 800 20472 79200 20872
rect 880 20192 79120 20472
rect 800 19656 79200 20192
rect 880 19376 79120 19656
rect 800 18840 79200 19376
rect 880 18560 79120 18840
rect 800 18024 79200 18560
rect 880 17744 79120 18024
rect 800 17208 79200 17744
rect 880 16928 79120 17208
rect 800 16392 79200 16928
rect 880 16112 79120 16392
rect 800 15576 79200 16112
rect 880 15296 79120 15576
rect 800 14760 79200 15296
rect 880 14480 79120 14760
rect 800 13944 79200 14480
rect 880 13664 79120 13944
rect 800 13264 79200 13664
rect 880 12984 79120 13264
rect 800 12448 79200 12984
rect 880 12168 79120 12448
rect 800 11632 79200 12168
rect 880 11352 79120 11632
rect 800 10816 79200 11352
rect 880 10536 79120 10816
rect 800 10000 79200 10536
rect 880 9720 79120 10000
rect 800 9184 79200 9720
rect 880 8904 79120 9184
rect 800 8368 79200 8904
rect 880 8088 79120 8368
rect 800 7552 79200 8088
rect 880 7272 79120 7552
rect 800 6872 79200 7272
rect 880 6592 79120 6872
rect 800 6056 79200 6592
rect 880 5776 79120 6056
rect 800 5240 79200 5776
rect 880 4960 79120 5240
rect 800 4424 79200 4960
rect 880 4144 79120 4424
rect 800 3608 79200 4144
rect 880 3328 79120 3608
rect 800 2792 79200 3328
rect 880 2512 79120 2792
rect 800 1976 79200 2512
rect 880 1696 79120 1976
rect 800 1160 79200 1696
rect 880 880 79120 1160
rect 800 480 79200 880
rect 880 307 79120 480
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< labels >>
rlabel metal2 s 78770 0 78826 800 6 io_wbs_ack
port 1 nsew signal output
rlabel metal3 s 79200 78616 80000 78736 6 io_wbs_ack_0
port 2 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 io_wbs_ack_1
port 3 nsew signal input
rlabel metal2 s 386 0 442 800 6 io_wbs_adr[0]
port 4 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_wbs_adr[10]
port 5 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 io_wbs_adr[11]
port 6 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 io_wbs_adr[12]
port 7 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 io_wbs_adr[13]
port 8 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 io_wbs_adr[14]
port 9 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 io_wbs_adr[15]
port 10 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 io_wbs_adr[16]
port 11 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 io_wbs_adr[17]
port 12 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 io_wbs_adr[18]
port 13 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 io_wbs_adr[19]
port 14 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 io_wbs_adr[1]
port 15 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 io_wbs_adr[20]
port 16 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 io_wbs_adr[21]
port 17 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 io_wbs_adr[22]
port 18 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 io_wbs_adr[23]
port 19 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 io_wbs_adr[24]
port 20 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 io_wbs_adr[25]
port 21 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 io_wbs_adr[26]
port 22 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_wbs_adr[27]
port 23 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 io_wbs_adr[28]
port 24 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 io_wbs_adr[29]
port 25 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 io_wbs_adr[2]
port 26 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 io_wbs_adr[30]
port 27 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 io_wbs_adr[31]
port 28 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 io_wbs_adr[3]
port 29 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 io_wbs_adr[4]
port 30 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 io_wbs_adr[5]
port 31 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_adr[6]
port 32 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 io_wbs_adr[7]
port 33 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 io_wbs_adr[8]
port 34 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 io_wbs_adr[9]
port 35 nsew signal input
rlabel metal3 s 79200 280 80000 400 6 io_wbs_adr_0[0]
port 36 nsew signal output
rlabel metal3 s 79200 8168 80000 8288 6 io_wbs_adr_0[10]
port 37 nsew signal output
rlabel metal3 s 79200 8984 80000 9104 6 io_wbs_adr_0[11]
port 38 nsew signal output
rlabel metal3 s 79200 9800 80000 9920 6 io_wbs_adr_0[12]
port 39 nsew signal output
rlabel metal3 s 79200 10616 80000 10736 6 io_wbs_adr_0[13]
port 40 nsew signal output
rlabel metal3 s 79200 11432 80000 11552 6 io_wbs_adr_0[14]
port 41 nsew signal output
rlabel metal3 s 79200 12248 80000 12368 6 io_wbs_adr_0[15]
port 42 nsew signal output
rlabel metal3 s 79200 13064 80000 13184 6 io_wbs_adr_0[16]
port 43 nsew signal output
rlabel metal3 s 79200 13744 80000 13864 6 io_wbs_adr_0[17]
port 44 nsew signal output
rlabel metal3 s 79200 14560 80000 14680 6 io_wbs_adr_0[18]
port 45 nsew signal output
rlabel metal3 s 79200 15376 80000 15496 6 io_wbs_adr_0[19]
port 46 nsew signal output
rlabel metal3 s 79200 960 80000 1080 6 io_wbs_adr_0[1]
port 47 nsew signal output
rlabel metal3 s 79200 16192 80000 16312 6 io_wbs_adr_0[20]
port 48 nsew signal output
rlabel metal3 s 79200 17008 80000 17128 6 io_wbs_adr_0[21]
port 49 nsew signal output
rlabel metal3 s 79200 17824 80000 17944 6 io_wbs_adr_0[22]
port 50 nsew signal output
rlabel metal3 s 79200 18640 80000 18760 6 io_wbs_adr_0[23]
port 51 nsew signal output
rlabel metal3 s 79200 19456 80000 19576 6 io_wbs_adr_0[24]
port 52 nsew signal output
rlabel metal3 s 79200 20272 80000 20392 6 io_wbs_adr_0[25]
port 53 nsew signal output
rlabel metal3 s 79200 20952 80000 21072 6 io_wbs_adr_0[26]
port 54 nsew signal output
rlabel metal3 s 79200 21768 80000 21888 6 io_wbs_adr_0[27]
port 55 nsew signal output
rlabel metal3 s 79200 22584 80000 22704 6 io_wbs_adr_0[28]
port 56 nsew signal output
rlabel metal3 s 79200 23400 80000 23520 6 io_wbs_adr_0[29]
port 57 nsew signal output
rlabel metal3 s 79200 1776 80000 1896 6 io_wbs_adr_0[2]
port 58 nsew signal output
rlabel metal3 s 79200 24216 80000 24336 6 io_wbs_adr_0[30]
port 59 nsew signal output
rlabel metal3 s 79200 25032 80000 25152 6 io_wbs_adr_0[31]
port 60 nsew signal output
rlabel metal3 s 79200 2592 80000 2712 6 io_wbs_adr_0[3]
port 61 nsew signal output
rlabel metal3 s 79200 3408 80000 3528 6 io_wbs_adr_0[4]
port 62 nsew signal output
rlabel metal3 s 79200 4224 80000 4344 6 io_wbs_adr_0[5]
port 63 nsew signal output
rlabel metal3 s 79200 5040 80000 5160 6 io_wbs_adr_0[6]
port 64 nsew signal output
rlabel metal3 s 79200 5856 80000 5976 6 io_wbs_adr_0[7]
port 65 nsew signal output
rlabel metal3 s 79200 6672 80000 6792 6 io_wbs_adr_0[8]
port 66 nsew signal output
rlabel metal3 s 79200 7352 80000 7472 6 io_wbs_adr_0[9]
port 67 nsew signal output
rlabel metal3 s 0 280 800 400 6 io_wbs_adr_1[0]
port 68 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_wbs_adr_1[10]
port 69 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 io_wbs_adr_1[11]
port 70 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_wbs_adr_1[12]
port 71 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 io_wbs_adr_1[13]
port 72 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 io_wbs_adr_1[14]
port 73 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_wbs_adr_1[15]
port 74 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 io_wbs_adr_1[16]
port 75 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 io_wbs_adr_1[17]
port 76 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 io_wbs_adr_1[18]
port 77 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 io_wbs_adr_1[19]
port 78 nsew signal output
rlabel metal3 s 0 960 800 1080 6 io_wbs_adr_1[1]
port 79 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 io_wbs_adr_1[20]
port 80 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 io_wbs_adr_1[21]
port 81 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 io_wbs_adr_1[22]
port 82 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 io_wbs_adr_1[23]
port 83 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 io_wbs_adr_1[24]
port 84 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 io_wbs_adr_1[25]
port 85 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 io_wbs_adr_1[26]
port 86 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_wbs_adr_1[27]
port 87 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 io_wbs_adr_1[28]
port 88 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_wbs_adr_1[29]
port 89 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_wbs_adr_1[2]
port 90 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 io_wbs_adr_1[30]
port 91 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 io_wbs_adr_1[31]
port 92 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 io_wbs_adr_1[3]
port 93 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 io_wbs_adr_1[4]
port 94 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_wbs_adr_1[5]
port 95 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 io_wbs_adr_1[6]
port 96 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 io_wbs_adr_1[7]
port 97 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_wbs_adr_1[8]
port 98 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 io_wbs_adr_1[9]
port 99 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 io_wbs_cyc
port 100 nsew signal input
rlabel metal3 s 79200 79432 80000 79552 6 io_wbs_cyc_0
port 101 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 io_wbs_cyc_1
port 102 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 io_wbs_datrd[0]
port 103 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 io_wbs_datrd[10]
port 104 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 io_wbs_datrd[11]
port 105 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 io_wbs_datrd[12]
port 106 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 io_wbs_datrd[13]
port 107 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 io_wbs_datrd[14]
port 108 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 io_wbs_datrd[15]
port 109 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_wbs_datrd[16]
port 110 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 io_wbs_datrd[17]
port 111 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 io_wbs_datrd[18]
port 112 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 io_wbs_datrd[19]
port 113 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 io_wbs_datrd[1]
port 114 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 io_wbs_datrd[20]
port 115 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 io_wbs_datrd[21]
port 116 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 io_wbs_datrd[22]
port 117 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 io_wbs_datrd[23]
port 118 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 io_wbs_datrd[24]
port 119 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 io_wbs_datrd[25]
port 120 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 io_wbs_datrd[26]
port 121 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 io_wbs_datrd[27]
port 122 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 io_wbs_datrd[28]
port 123 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 io_wbs_datrd[29]
port 124 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 io_wbs_datrd[2]
port 125 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 io_wbs_datrd[30]
port 126 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 io_wbs_datrd[31]
port 127 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 io_wbs_datrd[3]
port 128 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 io_wbs_datrd[4]
port 129 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 io_wbs_datrd[5]
port 130 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 io_wbs_datrd[6]
port 131 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 io_wbs_datrd[7]
port 132 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 io_wbs_datrd[8]
port 133 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 io_wbs_datrd[9]
port 134 nsew signal output
rlabel metal3 s 79200 51416 80000 51536 6 io_wbs_datrd_0[0]
port 135 nsew signal input
rlabel metal3 s 79200 59440 80000 59560 6 io_wbs_datrd_0[10]
port 136 nsew signal input
rlabel metal3 s 79200 60256 80000 60376 6 io_wbs_datrd_0[11]
port 137 nsew signal input
rlabel metal3 s 79200 60936 80000 61056 6 io_wbs_datrd_0[12]
port 138 nsew signal input
rlabel metal3 s 79200 61752 80000 61872 6 io_wbs_datrd_0[13]
port 139 nsew signal input
rlabel metal3 s 79200 62568 80000 62688 6 io_wbs_datrd_0[14]
port 140 nsew signal input
rlabel metal3 s 79200 63384 80000 63504 6 io_wbs_datrd_0[15]
port 141 nsew signal input
rlabel metal3 s 79200 64200 80000 64320 6 io_wbs_datrd_0[16]
port 142 nsew signal input
rlabel metal3 s 79200 65016 80000 65136 6 io_wbs_datrd_0[17]
port 143 nsew signal input
rlabel metal3 s 79200 65832 80000 65952 6 io_wbs_datrd_0[18]
port 144 nsew signal input
rlabel metal3 s 79200 66648 80000 66768 6 io_wbs_datrd_0[19]
port 145 nsew signal input
rlabel metal3 s 79200 52232 80000 52352 6 io_wbs_datrd_0[1]
port 146 nsew signal input
rlabel metal3 s 79200 67328 80000 67448 6 io_wbs_datrd_0[20]
port 147 nsew signal input
rlabel metal3 s 79200 68144 80000 68264 6 io_wbs_datrd_0[21]
port 148 nsew signal input
rlabel metal3 s 79200 68960 80000 69080 6 io_wbs_datrd_0[22]
port 149 nsew signal input
rlabel metal3 s 79200 69776 80000 69896 6 io_wbs_datrd_0[23]
port 150 nsew signal input
rlabel metal3 s 79200 70592 80000 70712 6 io_wbs_datrd_0[24]
port 151 nsew signal input
rlabel metal3 s 79200 71408 80000 71528 6 io_wbs_datrd_0[25]
port 152 nsew signal input
rlabel metal3 s 79200 72224 80000 72344 6 io_wbs_datrd_0[26]
port 153 nsew signal input
rlabel metal3 s 79200 73040 80000 73160 6 io_wbs_datrd_0[27]
port 154 nsew signal input
rlabel metal3 s 79200 73720 80000 73840 6 io_wbs_datrd_0[28]
port 155 nsew signal input
rlabel metal3 s 79200 74536 80000 74656 6 io_wbs_datrd_0[29]
port 156 nsew signal input
rlabel metal3 s 79200 53048 80000 53168 6 io_wbs_datrd_0[2]
port 157 nsew signal input
rlabel metal3 s 79200 75352 80000 75472 6 io_wbs_datrd_0[30]
port 158 nsew signal input
rlabel metal3 s 79200 76168 80000 76288 6 io_wbs_datrd_0[31]
port 159 nsew signal input
rlabel metal3 s 79200 53728 80000 53848 6 io_wbs_datrd_0[3]
port 160 nsew signal input
rlabel metal3 s 79200 54544 80000 54664 6 io_wbs_datrd_0[4]
port 161 nsew signal input
rlabel metal3 s 79200 55360 80000 55480 6 io_wbs_datrd_0[5]
port 162 nsew signal input
rlabel metal3 s 79200 56176 80000 56296 6 io_wbs_datrd_0[6]
port 163 nsew signal input
rlabel metal3 s 79200 56992 80000 57112 6 io_wbs_datrd_0[7]
port 164 nsew signal input
rlabel metal3 s 79200 57808 80000 57928 6 io_wbs_datrd_0[8]
port 165 nsew signal input
rlabel metal3 s 79200 58624 80000 58744 6 io_wbs_datrd_0[9]
port 166 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 io_wbs_datrd_1[0]
port 167 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 io_wbs_datrd_1[10]
port 168 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 io_wbs_datrd_1[11]
port 169 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 io_wbs_datrd_1[12]
port 170 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 io_wbs_datrd_1[13]
port 171 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 io_wbs_datrd_1[14]
port 172 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 io_wbs_datrd_1[15]
port 173 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 io_wbs_datrd_1[16]
port 174 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 io_wbs_datrd_1[17]
port 175 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 io_wbs_datrd_1[18]
port 176 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 io_wbs_datrd_1[19]
port 177 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 io_wbs_datrd_1[1]
port 178 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 io_wbs_datrd_1[20]
port 179 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 io_wbs_datrd_1[21]
port 180 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 io_wbs_datrd_1[22]
port 181 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 io_wbs_datrd_1[23]
port 182 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 io_wbs_datrd_1[24]
port 183 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 io_wbs_datrd_1[25]
port 184 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 io_wbs_datrd_1[26]
port 185 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 io_wbs_datrd_1[27]
port 186 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 io_wbs_datrd_1[28]
port 187 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 io_wbs_datrd_1[29]
port 188 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_wbs_datrd_1[2]
port 189 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 io_wbs_datrd_1[30]
port 190 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 io_wbs_datrd_1[31]
port 191 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 io_wbs_datrd_1[3]
port 192 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 io_wbs_datrd_1[4]
port 193 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 io_wbs_datrd_1[5]
port 194 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 io_wbs_datrd_1[6]
port 195 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 io_wbs_datrd_1[7]
port 196 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 io_wbs_datrd_1[8]
port 197 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 io_wbs_datrd_1[9]
port 198 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 io_wbs_datwr[0]
port 199 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 io_wbs_datwr[10]
port 200 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 io_wbs_datwr[11]
port 201 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 io_wbs_datwr[12]
port 202 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 io_wbs_datwr[13]
port 203 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 io_wbs_datwr[14]
port 204 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 io_wbs_datwr[15]
port 205 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 io_wbs_datwr[16]
port 206 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 io_wbs_datwr[17]
port 207 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 io_wbs_datwr[18]
port 208 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 io_wbs_datwr[19]
port 209 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 io_wbs_datwr[1]
port 210 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 io_wbs_datwr[20]
port 211 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 io_wbs_datwr[21]
port 212 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 io_wbs_datwr[22]
port 213 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 io_wbs_datwr[23]
port 214 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 io_wbs_datwr[24]
port 215 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 io_wbs_datwr[25]
port 216 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 io_wbs_datwr[26]
port 217 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 io_wbs_datwr[27]
port 218 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 io_wbs_datwr[28]
port 219 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 io_wbs_datwr[29]
port 220 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 io_wbs_datwr[2]
port 221 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 io_wbs_datwr[30]
port 222 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 io_wbs_datwr[31]
port 223 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_wbs_datwr[3]
port 224 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 io_wbs_datwr[4]
port 225 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 io_wbs_datwr[5]
port 226 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 io_wbs_datwr[6]
port 227 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 io_wbs_datwr[7]
port 228 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 io_wbs_datwr[8]
port 229 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 io_wbs_datwr[9]
port 230 nsew signal input
rlabel metal3 s 79200 25848 80000 25968 6 io_wbs_datwr_0[0]
port 231 nsew signal output
rlabel metal3 s 79200 33736 80000 33856 6 io_wbs_datwr_0[10]
port 232 nsew signal output
rlabel metal3 s 79200 34552 80000 34672 6 io_wbs_datwr_0[11]
port 233 nsew signal output
rlabel metal3 s 79200 35368 80000 35488 6 io_wbs_datwr_0[12]
port 234 nsew signal output
rlabel metal3 s 79200 36184 80000 36304 6 io_wbs_datwr_0[13]
port 235 nsew signal output
rlabel metal3 s 79200 37000 80000 37120 6 io_wbs_datwr_0[14]
port 236 nsew signal output
rlabel metal3 s 79200 37816 80000 37936 6 io_wbs_datwr_0[15]
port 237 nsew signal output
rlabel metal3 s 79200 38632 80000 38752 6 io_wbs_datwr_0[16]
port 238 nsew signal output
rlabel metal3 s 79200 39448 80000 39568 6 io_wbs_datwr_0[17]
port 239 nsew signal output
rlabel metal3 s 79200 40264 80000 40384 6 io_wbs_datwr_0[18]
port 240 nsew signal output
rlabel metal3 s 79200 40944 80000 41064 6 io_wbs_datwr_0[19]
port 241 nsew signal output
rlabel metal3 s 79200 26664 80000 26784 6 io_wbs_datwr_0[1]
port 242 nsew signal output
rlabel metal3 s 79200 41760 80000 41880 6 io_wbs_datwr_0[20]
port 243 nsew signal output
rlabel metal3 s 79200 42576 80000 42696 6 io_wbs_datwr_0[21]
port 244 nsew signal output
rlabel metal3 s 79200 43392 80000 43512 6 io_wbs_datwr_0[22]
port 245 nsew signal output
rlabel metal3 s 79200 44208 80000 44328 6 io_wbs_datwr_0[23]
port 246 nsew signal output
rlabel metal3 s 79200 45024 80000 45144 6 io_wbs_datwr_0[24]
port 247 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 io_wbs_datwr_0[25]
port 248 nsew signal output
rlabel metal3 s 79200 46656 80000 46776 6 io_wbs_datwr_0[26]
port 249 nsew signal output
rlabel metal3 s 79200 47336 80000 47456 6 io_wbs_datwr_0[27]
port 250 nsew signal output
rlabel metal3 s 79200 48152 80000 48272 6 io_wbs_datwr_0[28]
port 251 nsew signal output
rlabel metal3 s 79200 48968 80000 49088 6 io_wbs_datwr_0[29]
port 252 nsew signal output
rlabel metal3 s 79200 27344 80000 27464 6 io_wbs_datwr_0[2]
port 253 nsew signal output
rlabel metal3 s 79200 49784 80000 49904 6 io_wbs_datwr_0[30]
port 254 nsew signal output
rlabel metal3 s 79200 50600 80000 50720 6 io_wbs_datwr_0[31]
port 255 nsew signal output
rlabel metal3 s 79200 28160 80000 28280 6 io_wbs_datwr_0[3]
port 256 nsew signal output
rlabel metal3 s 79200 28976 80000 29096 6 io_wbs_datwr_0[4]
port 257 nsew signal output
rlabel metal3 s 79200 29792 80000 29912 6 io_wbs_datwr_0[5]
port 258 nsew signal output
rlabel metal3 s 79200 30608 80000 30728 6 io_wbs_datwr_0[6]
port 259 nsew signal output
rlabel metal3 s 79200 31424 80000 31544 6 io_wbs_datwr_0[7]
port 260 nsew signal output
rlabel metal3 s 79200 32240 80000 32360 6 io_wbs_datwr_0[8]
port 261 nsew signal output
rlabel metal3 s 79200 33056 80000 33176 6 io_wbs_datwr_0[9]
port 262 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_wbs_datwr_1[0]
port 263 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 io_wbs_datwr_1[10]
port 264 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 io_wbs_datwr_1[11]
port 265 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_wbs_datwr_1[12]
port 266 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 io_wbs_datwr_1[13]
port 267 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 io_wbs_datwr_1[14]
port 268 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 io_wbs_datwr_1[15]
port 269 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 io_wbs_datwr_1[16]
port 270 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_wbs_datwr_1[17]
port 271 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 io_wbs_datwr_1[18]
port 272 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 io_wbs_datwr_1[19]
port 273 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_wbs_datwr_1[1]
port 274 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 io_wbs_datwr_1[20]
port 275 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 io_wbs_datwr_1[21]
port 276 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_wbs_datwr_1[22]
port 277 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_wbs_datwr_1[23]
port 278 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 io_wbs_datwr_1[24]
port 279 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_wbs_datwr_1[25]
port 280 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 io_wbs_datwr_1[26]
port 281 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_wbs_datwr_1[27]
port 282 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 io_wbs_datwr_1[28]
port 283 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 io_wbs_datwr_1[29]
port 284 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 io_wbs_datwr_1[2]
port 285 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 io_wbs_datwr_1[30]
port 286 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 io_wbs_datwr_1[31]
port 287 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 io_wbs_datwr_1[3]
port 288 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 io_wbs_datwr_1[4]
port 289 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 io_wbs_datwr_1[5]
port 290 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 io_wbs_datwr_1[6]
port 291 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 io_wbs_datwr_1[7]
port 292 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 io_wbs_datwr_1[8]
port 293 nsew signal output
rlabel metal3 s 0 33056 800 33176 6 io_wbs_datwr_1[9]
port 294 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 io_wbs_stb
port 295 nsew signal input
rlabel metal3 s 79200 77800 80000 77920 6 io_wbs_stb_0
port 296 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 io_wbs_stb_1
port 297 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 io_wbs_we
port 298 nsew signal input
rlabel metal3 s 79200 76984 80000 77104 6 io_wbs_we_0
port 299 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 io_wbs_we_1
port 300 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 301 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 301 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 301 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 302 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 302 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2731750
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/wb_mux/runs/wb_mux/results/finishing/wb_mux.magic.gds
string GDS_START 115078
<< end >>

