magic
tech sky130A
magscale 1 2
timestamp 1657200204
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 407114 700408 407120 700460
rect 407172 700448 407178 700460
rect 478506 700448 478512 700460
rect 407172 700420 478512 700448
rect 407172 700408 407178 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 517514 700408 517520 700460
rect 517572 700448 517578 700460
rect 527174 700448 527180 700460
rect 517572 700420 527180 700448
rect 517572 700408 517578 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 397454 700340 397460 700392
rect 397512 700380 397518 700392
rect 524414 700380 524420 700392
rect 397512 700352 524420 700380
rect 397512 700340 397518 700352
rect 524414 700340 524420 700352
rect 524472 700340 524478 700392
rect 404354 700272 404360 700324
rect 404412 700312 404418 700324
rect 543458 700312 543464 700324
rect 404412 700284 543464 700312
rect 404412 700272 404418 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 409874 699660 409880 699712
rect 409932 699700 409938 699712
rect 413646 699700 413652 699712
rect 409932 699672 413652 699700
rect 409932 699660 409938 699672
rect 413646 699660 413652 699672
rect 413704 699660 413710 699712
rect 514754 696940 514760 696992
rect 514812 696980 514818 696992
rect 580166 696980 580172 696992
rect 514812 696952 580172 696980
rect 514812 696940 514818 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 400214 683136 400220 683188
rect 400272 683176 400278 683188
rect 580166 683176 580172 683188
rect 400272 683148 580172 683176
rect 400272 683136 400278 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 510614 643084 510620 643136
rect 510672 643124 510678 643136
rect 580166 643124 580172 643136
rect 510672 643096 580172 643124
rect 510672 643084 510678 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 397454 630640 397460 630692
rect 397512 630680 397518 630692
rect 580166 630680 580172 630692
rect 397512 630652 580172 630680
rect 397512 630640 397518 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 507854 590656 507860 590708
rect 507912 590696 507918 590708
rect 579798 590696 579804 590708
rect 507912 590668 579804 590696
rect 507912 590656 507918 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 393314 576852 393320 576904
rect 393372 576892 393378 576904
rect 580166 576892 580172 576904
rect 393372 576864 580172 576892
rect 393372 576852 393378 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 347774 552712 347780 552764
rect 347832 552752 347838 552764
rect 414014 552752 414020 552764
rect 347832 552724 414020 552752
rect 347832 552712 347838 552724
rect 414014 552712 414020 552724
rect 414072 552712 414078 552764
rect 462314 552712 462320 552764
rect 462372 552752 462378 552764
rect 521654 552752 521660 552764
rect 462372 552724 521660 552752
rect 462372 552712 462378 552724
rect 521654 552712 521660 552724
rect 521712 552712 521718 552764
rect 331214 552644 331220 552696
rect 331272 552684 331278 552696
rect 527910 552684 527916 552696
rect 331272 552656 527916 552684
rect 331272 552644 331278 552656
rect 527910 552644 527916 552656
rect 527968 552644 527974 552696
rect 505738 552440 505744 552492
rect 505796 552480 505802 552492
rect 547138 552480 547144 552492
rect 505796 552452 547144 552480
rect 505796 552440 505802 552452
rect 547138 552440 547144 552452
rect 547196 552440 547202 552492
rect 499206 552372 499212 552424
rect 499264 552412 499270 552424
rect 551278 552412 551284 552424
rect 499264 552384 551284 552412
rect 499264 552372 499270 552384
rect 551278 552372 551284 552384
rect 551336 552372 551342 552424
rect 495986 552304 495992 552356
rect 496044 552344 496050 552356
rect 548518 552344 548524 552356
rect 496044 552316 548524 552344
rect 496044 552304 496050 552316
rect 548518 552304 548524 552316
rect 548576 552304 548582 552356
rect 391658 552236 391664 552288
rect 391716 552276 391722 552288
rect 555418 552276 555424 552288
rect 391716 552248 555424 552276
rect 391716 552236 391722 552248
rect 555418 552236 555424 552248
rect 555476 552236 555482 552288
rect 388346 552168 388352 552220
rect 388404 552208 388410 552220
rect 554038 552208 554044 552220
rect 388404 552180 554044 552208
rect 388404 552168 388410 552180
rect 554038 552168 554044 552180
rect 554096 552168 554102 552220
rect 384942 552100 384948 552152
rect 385000 552140 385006 552152
rect 556798 552140 556804 552152
rect 385000 552112 556804 552140
rect 385000 552100 385006 552112
rect 556798 552100 556804 552112
rect 556856 552100 556862 552152
rect 381906 552032 381912 552084
rect 381964 552072 381970 552084
rect 558178 552072 558184 552084
rect 381964 552044 558184 552072
rect 381964 552032 381970 552044
rect 558178 552032 558184 552044
rect 558236 552032 558242 552084
rect 502334 549244 502340 549296
rect 502392 549284 502398 549296
rect 580258 549284 580264 549296
rect 502392 549256 580264 549284
rect 502392 549244 502398 549256
rect 580258 549244 580264 549256
rect 580316 549244 580322 549296
rect 268378 547884 268384 547936
rect 268436 547924 268442 547936
rect 376938 547924 376944 547936
rect 268436 547896 376944 547924
rect 268436 547884 268442 547896
rect 376938 547884 376944 547896
rect 376996 547884 377002 547936
rect 251818 545096 251824 545148
rect 251876 545136 251882 545148
rect 376938 545136 376944 545148
rect 251876 545108 376944 545136
rect 251876 545096 251882 545108
rect 376938 545096 376944 545108
rect 376996 545096 377002 545148
rect 266998 542376 267004 542428
rect 267056 542416 267062 542428
rect 376846 542416 376852 542428
rect 267056 542388 376852 542416
rect 267056 542376 267062 542388
rect 376846 542376 376852 542388
rect 376904 542376 376910 542428
rect 264238 538228 264244 538280
rect 264296 538268 264302 538280
rect 376938 538268 376944 538280
rect 264296 538240 376944 538268
rect 264296 538228 264302 538240
rect 376938 538228 376944 538240
rect 376996 538228 377002 538280
rect 547138 538160 547144 538212
rect 547196 538200 547202 538212
rect 579890 538200 579896 538212
rect 547196 538172 579896 538200
rect 547196 538160 547202 538172
rect 579890 538160 579896 538172
rect 579948 538160 579954 538212
rect 251910 535440 251916 535492
rect 251968 535480 251974 535492
rect 376938 535480 376944 535492
rect 251968 535452 376944 535480
rect 251968 535440 251974 535452
rect 376938 535440 376944 535452
rect 376996 535440 377002 535492
rect 262858 532720 262864 532772
rect 262916 532760 262922 532772
rect 376938 532760 376944 532772
rect 262916 532732 376944 532760
rect 262916 532720 262922 532732
rect 376938 532720 376944 532732
rect 376996 532720 377002 532772
rect 260098 527144 260104 527196
rect 260156 527184 260162 527196
rect 376938 527184 376944 527196
rect 260156 527156 376944 527184
rect 260156 527144 260162 527156
rect 376938 527144 376944 527156
rect 376996 527144 377002 527196
rect 555418 525716 555424 525768
rect 555476 525756 555482 525768
rect 580166 525756 580172 525768
rect 555476 525728 580172 525756
rect 555476 525716 555482 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 252002 524424 252008 524476
rect 252060 524464 252066 524476
rect 376938 524464 376944 524476
rect 252060 524436 376944 524464
rect 252060 524424 252066 524436
rect 376938 524424 376944 524436
rect 376996 524424 377002 524476
rect 258718 522996 258724 523048
rect 258776 523036 258782 523048
rect 376938 523036 376944 523048
rect 258776 523008 376944 523036
rect 258776 522996 258782 523008
rect 376938 522996 376944 523008
rect 376996 522996 377002 523048
rect 255958 517488 255964 517540
rect 256016 517528 256022 517540
rect 376938 517528 376944 517540
rect 256016 517500 376944 517528
rect 256016 517488 256022 517500
rect 376938 517488 376944 517500
rect 376996 517488 377002 517540
rect 252094 514768 252100 514820
rect 252152 514808 252158 514820
rect 376938 514808 376944 514820
rect 252152 514780 376944 514808
rect 252152 514768 252158 514780
rect 376938 514768 376944 514780
rect 376996 514768 377002 514820
rect 253198 511980 253204 512032
rect 253256 512020 253262 512032
rect 376938 512020 376944 512032
rect 253256 511992 376944 512020
rect 253256 511980 253262 511992
rect 376938 511980 376944 511992
rect 376996 511980 377002 512032
rect 253290 509260 253296 509312
rect 253348 509300 253354 509312
rect 376938 509300 376944 509312
rect 253348 509272 376944 509300
rect 253348 509260 253354 509272
rect 376938 509260 376944 509272
rect 376996 509260 377002 509312
rect 252462 499468 252468 499520
rect 252520 499508 252526 499520
rect 268378 499508 268384 499520
rect 252520 499480 268384 499508
rect 252520 499468 252526 499480
rect 268378 499468 268384 499480
rect 268436 499468 268442 499520
rect 252462 498108 252468 498160
rect 252520 498148 252526 498160
rect 266998 498148 267004 498160
rect 252520 498120 267004 498148
rect 252520 498108 252526 498120
rect 266998 498108 267004 498120
rect 267056 498108 267062 498160
rect 252462 496748 252468 496800
rect 252520 496788 252526 496800
rect 377398 496788 377404 496800
rect 252520 496760 377404 496788
rect 252520 496748 252526 496760
rect 377398 496748 377404 496760
rect 377456 496748 377462 496800
rect 252370 496680 252376 496732
rect 252428 496720 252434 496732
rect 264238 496720 264244 496732
rect 252428 496692 264244 496720
rect 252428 496680 252434 496692
rect 264238 496680 264244 496692
rect 264296 496680 264302 496732
rect 377306 494708 377312 494760
rect 377364 494748 377370 494760
rect 377766 494748 377772 494760
rect 377364 494720 377772 494748
rect 377364 494708 377370 494720
rect 377766 494708 377772 494720
rect 377824 494708 377830 494760
rect 252370 493960 252376 494012
rect 252428 494000 252434 494012
rect 377490 494000 377496 494012
rect 252428 493972 377496 494000
rect 252428 493960 252434 493972
rect 377490 493960 377496 493972
rect 377548 493960 377554 494012
rect 252462 493892 252468 493944
rect 252520 493932 252526 493944
rect 262858 493932 262864 493944
rect 252520 493904 262864 493932
rect 252520 493892 252526 493904
rect 262858 493892 262864 493904
rect 262916 493892 262922 493944
rect 252462 491988 252468 492040
rect 252520 492028 252526 492040
rect 260098 492028 260104 492040
rect 252520 492000 260104 492028
rect 252520 491988 252526 492000
rect 260098 491988 260104 492000
rect 260156 491988 260162 492040
rect 251818 491308 251824 491360
rect 251876 491348 251882 491360
rect 376938 491348 376944 491360
rect 251876 491320 376944 491348
rect 251876 491308 251882 491320
rect 376938 491308 376944 491320
rect 376996 491308 377002 491360
rect 251910 491172 251916 491224
rect 251968 491212 251974 491224
rect 258718 491212 258724 491224
rect 251968 491184 258724 491212
rect 251968 491172 251974 491184
rect 258718 491172 258724 491184
rect 258776 491172 258782 491224
rect 252462 489812 252468 489864
rect 252520 489852 252526 489864
rect 377582 489852 377588 489864
rect 252520 489824 377588 489852
rect 252520 489812 252526 489824
rect 377582 489812 377588 489824
rect 377640 489812 377646 489864
rect 252002 488520 252008 488572
rect 252060 488560 252066 488572
rect 376938 488560 376944 488572
rect 252060 488532 376944 488560
rect 252060 488520 252066 488532
rect 376938 488520 376944 488532
rect 376996 488520 377002 488572
rect 252462 488452 252468 488504
rect 252520 488492 252526 488504
rect 255958 488492 255964 488504
rect 252520 488464 255964 488492
rect 252520 488452 252526 488464
rect 255958 488452 255964 488464
rect 256016 488452 256022 488504
rect 251910 487160 251916 487212
rect 251968 487200 251974 487212
rect 376938 487200 376944 487212
rect 251968 487172 376944 487200
rect 251968 487160 251974 487172
rect 376938 487160 376944 487172
rect 376996 487160 377002 487212
rect 251266 487092 251272 487144
rect 251324 487132 251330 487144
rect 253198 487132 253204 487144
rect 251324 487104 253204 487132
rect 251324 487092 251330 487104
rect 253198 487092 253204 487104
rect 253256 487092 253262 487144
rect 251726 485732 251732 485784
rect 251784 485772 251790 485784
rect 377674 485772 377680 485784
rect 251784 485744 377680 485772
rect 251784 485732 251790 485744
rect 377674 485732 377680 485744
rect 377732 485732 377738 485784
rect 251358 485596 251364 485648
rect 251416 485636 251422 485648
rect 253290 485636 253296 485648
rect 251416 485608 253296 485636
rect 251416 485596 251422 485608
rect 253290 485596 253296 485608
rect 253348 485596 253354 485648
rect 251726 484304 251732 484356
rect 251784 484344 251790 484356
rect 377306 484344 377312 484356
rect 251784 484316 377312 484344
rect 251784 484304 251790 484316
rect 377306 484304 377312 484316
rect 377364 484304 377370 484356
rect 252462 482944 252468 482996
rect 252520 482984 252526 482996
rect 377858 482984 377864 482996
rect 252520 482956 377864 482984
rect 252520 482944 252526 482956
rect 377858 482944 377864 482956
rect 377916 482944 377922 482996
rect 252370 482876 252376 482928
rect 252428 482916 252434 482928
rect 377950 482916 377956 482928
rect 252428 482888 377956 482916
rect 252428 482876 252434 482888
rect 377950 482876 377956 482888
rect 378008 482876 378014 482928
rect 251726 481584 251732 481636
rect 251784 481624 251790 481636
rect 378042 481624 378048 481636
rect 251784 481596 378048 481624
rect 251784 481584 251790 481596
rect 378042 481584 378048 481596
rect 378100 481584 378106 481636
rect 252462 480156 252468 480208
rect 252520 480196 252526 480208
rect 377398 480196 377404 480208
rect 252520 480168 377404 480196
rect 252520 480156 252526 480168
rect 377398 480156 377404 480168
rect 377456 480156 377462 480208
rect 251726 477436 251732 477488
rect 251784 477476 251790 477488
rect 377490 477476 377496 477488
rect 251784 477448 377496 477476
rect 251784 477436 251790 477448
rect 377490 477436 377496 477448
rect 377548 477436 377554 477488
rect 251910 476076 251916 476128
rect 251968 476116 251974 476128
rect 376938 476116 376944 476128
rect 251968 476088 376944 476116
rect 251968 476076 251974 476088
rect 376938 476076 376944 476088
rect 376996 476076 377002 476128
rect 252462 476008 252468 476060
rect 252520 476048 252526 476060
rect 377214 476048 377220 476060
rect 252520 476020 377220 476048
rect 252520 476008 252526 476020
rect 377214 476008 377220 476020
rect 377272 476008 377278 476060
rect 252462 474648 252468 474700
rect 252520 474688 252526 474700
rect 377030 474688 377036 474700
rect 252520 474660 377036 474688
rect 252520 474648 252526 474660
rect 377030 474648 377036 474660
rect 377088 474648 377094 474700
rect 251542 473356 251548 473408
rect 251600 473396 251606 473408
rect 376938 473396 376944 473408
rect 251600 473368 376944 473396
rect 251600 473356 251606 473368
rect 376938 473356 376944 473368
rect 376996 473356 377002 473408
rect 554038 471928 554044 471980
rect 554096 471968 554102 471980
rect 580166 471968 580172 471980
rect 554096 471940 580172 471968
rect 554096 471928 554102 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 252462 471248 252468 471300
rect 252520 471288 252526 471300
rect 376938 471288 376944 471300
rect 252520 471260 376944 471288
rect 252520 471248 252526 471260
rect 376938 471248 376944 471260
rect 376996 471248 377002 471300
rect 252462 470500 252468 470552
rect 252520 470540 252526 470552
rect 376938 470540 376944 470552
rect 252520 470512 376944 470540
rect 252520 470500 252526 470512
rect 376938 470500 376944 470512
rect 376996 470500 377002 470552
rect 252462 467780 252468 467832
rect 252520 467820 252526 467832
rect 376938 467820 376944 467832
rect 252520 467792 376944 467820
rect 252520 467780 252526 467792
rect 376938 467780 376944 467792
rect 376996 467780 377002 467832
rect 252370 464992 252376 465044
rect 252428 465032 252434 465044
rect 376938 465032 376944 465044
rect 252428 465004 376944 465032
rect 252428 464992 252434 465004
rect 376938 464992 376944 465004
rect 376996 464992 377002 465044
rect 251266 463768 251272 463820
rect 251324 463808 251330 463820
rect 253198 463808 253204 463820
rect 251324 463780 253204 463808
rect 251324 463768 251330 463780
rect 253198 463768 253204 463780
rect 253256 463768 253262 463820
rect 251542 462272 251548 462324
rect 251600 462312 251606 462324
rect 376938 462312 376944 462324
rect 251600 462284 376944 462312
rect 251600 462272 251606 462284
rect 376938 462272 376944 462284
rect 376996 462272 377002 462324
rect 252462 459484 252468 459536
rect 252520 459524 252526 459536
rect 376938 459524 376944 459536
rect 252520 459496 376944 459524
rect 252520 459484 252526 459496
rect 376938 459484 376944 459496
rect 376996 459484 377002 459536
rect 143442 458056 143448 458108
rect 143500 458096 143506 458108
rect 218698 458096 218704 458108
rect 143500 458068 218704 458096
rect 143500 458056 143506 458068
rect 218698 458056 218704 458068
rect 218756 458056 218762 458108
rect 142062 457988 142068 458040
rect 142120 458028 142126 458040
rect 218790 458028 218796 458040
rect 142120 458000 218796 458028
rect 142120 457988 142126 458000
rect 218790 457988 218796 458000
rect 218848 457988 218854 458040
rect 152458 457920 152464 457972
rect 152516 457960 152522 457972
rect 239122 457960 239128 457972
rect 152516 457932 239128 457960
rect 152516 457920 152522 457932
rect 239122 457920 239128 457932
rect 239180 457920 239186 457972
rect 155218 457852 155224 457904
rect 155276 457892 155282 457904
rect 249150 457892 249156 457904
rect 155276 457864 249156 457892
rect 155276 457852 155282 457864
rect 249150 457852 249156 457864
rect 249208 457852 249214 457904
rect 140038 457784 140044 457836
rect 140096 457824 140102 457836
rect 244826 457824 244832 457836
rect 140096 457796 244832 457824
rect 140096 457784 140102 457796
rect 244826 457784 244832 457796
rect 244884 457784 244890 457836
rect 134518 457716 134524 457768
rect 134576 457756 134582 457768
rect 241974 457756 241980 457768
rect 134576 457728 241980 457756
rect 134576 457716 134582 457728
rect 241974 457716 241980 457728
rect 242032 457716 242038 457768
rect 90358 457648 90364 457700
rect 90416 457688 90422 457700
rect 216306 457688 216312 457700
rect 90416 457660 216312 457688
rect 90416 457648 90422 457660
rect 216306 457648 216312 457660
rect 216364 457648 216370 457700
rect 86218 457580 86224 457632
rect 86276 457620 86282 457632
rect 213454 457620 213460 457632
rect 86276 457592 213460 457620
rect 86276 457580 86282 457592
rect 213454 457580 213460 457592
rect 213512 457580 213518 457632
rect 79318 457512 79324 457564
rect 79376 457552 79382 457564
rect 207750 457552 207756 457564
rect 79376 457524 207756 457552
rect 79376 457512 79382 457524
rect 207750 457512 207756 457524
rect 207808 457512 207814 457564
rect 218882 457512 218888 457564
rect 218940 457552 218946 457564
rect 240594 457552 240600 457564
rect 218940 457524 240600 457552
rect 218940 457512 218946 457524
rect 240594 457512 240600 457524
rect 240652 457512 240658 457564
rect 80698 457444 80704 457496
rect 80756 457484 80762 457496
rect 210602 457484 210608 457496
rect 80756 457456 210608 457484
rect 80756 457444 80762 457456
rect 210602 457444 210608 457456
rect 210660 457444 210666 457496
rect 220078 457444 220084 457496
rect 220136 457484 220142 457496
rect 243446 457484 243452 457496
rect 220136 457456 243452 457484
rect 220136 457444 220142 457456
rect 243446 457444 243452 457456
rect 243504 457444 243510 457496
rect 252278 456696 252284 456748
rect 252336 456736 252342 456748
rect 376938 456736 376944 456748
rect 252336 456708 376944 456736
rect 252336 456696 252342 456708
rect 376938 456696 376944 456708
rect 376996 456696 377002 456748
rect 253198 455336 253204 455388
rect 253256 455376 253262 455388
rect 376938 455376 376944 455388
rect 253256 455348 376944 455376
rect 253256 455336 253262 455348
rect 376938 455336 376944 455348
rect 376996 455336 377002 455388
rect 252186 452548 252192 452600
rect 252244 452588 252250 452600
rect 376846 452588 376852 452600
rect 252244 452560 376852 452588
rect 252244 452548 252250 452560
rect 376846 452548 376852 452560
rect 376904 452548 376910 452600
rect 252002 449828 252008 449880
rect 252060 449868 252066 449880
rect 376938 449868 376944 449880
rect 252060 449840 376944 449868
rect 252060 449828 252066 449840
rect 376938 449828 376944 449840
rect 376996 449828 377002 449880
rect 252094 447040 252100 447092
rect 252152 447080 252158 447092
rect 376938 447080 376944 447092
rect 252152 447052 376944 447080
rect 252152 447040 252158 447052
rect 376938 447040 376944 447052
rect 376996 447040 377002 447092
rect 251910 444320 251916 444372
rect 251968 444360 251974 444372
rect 376846 444360 376852 444372
rect 251968 444332 376852 444360
rect 251968 444320 251974 444332
rect 376846 444320 376852 444332
rect 376904 444320 376910 444372
rect 251818 441532 251824 441584
rect 251876 441572 251882 441584
rect 376938 441572 376944 441584
rect 251876 441544 376944 441572
rect 251876 441532 251882 441544
rect 376938 441532 376944 441544
rect 376996 441532 377002 441584
rect 465718 438676 465724 438728
rect 465776 438716 465782 438728
rect 498194 438716 498200 438728
rect 465776 438688 498200 438716
rect 465776 438676 465782 438688
rect 498194 438676 498200 438688
rect 498252 438676 498258 438728
rect 461578 438608 461584 438660
rect 461636 438648 461642 438660
rect 480346 438648 480352 438660
rect 461636 438620 480352 438648
rect 461636 438608 461642 438620
rect 480346 438608 480352 438620
rect 480404 438608 480410 438660
rect 482278 438608 482284 438660
rect 482336 438648 482342 438660
rect 525886 438648 525892 438660
rect 482336 438620 525892 438648
rect 482336 438608 482342 438620
rect 525886 438608 525892 438620
rect 525944 438608 525950 438660
rect 395338 438540 395344 438592
rect 395396 438580 395402 438592
rect 408494 438580 408500 438592
rect 395396 438552 408500 438580
rect 395396 438540 395402 438552
rect 408494 438540 408500 438552
rect 408552 438540 408558 438592
rect 468478 438540 468484 438592
rect 468536 438580 468542 438592
rect 512638 438580 512644 438592
rect 468536 438552 512644 438580
rect 468536 438540 468542 438552
rect 512638 438540 512644 438552
rect 512696 438540 512702 438592
rect 381538 438472 381544 438524
rect 381596 438512 381602 438524
rect 397914 438512 397920 438524
rect 381596 438484 397920 438512
rect 381596 438472 381602 438484
rect 397914 438472 397920 438484
rect 397972 438472 397978 438524
rect 453298 438472 453304 438524
rect 453356 438512 453362 438524
rect 462590 438512 462596 438524
rect 453356 438484 462596 438512
rect 453356 438472 453362 438484
rect 462590 438472 462596 438484
rect 462648 438472 462654 438524
rect 464338 438472 464344 438524
rect 464396 438512 464402 438524
rect 508222 438512 508228 438524
rect 464396 438484 508228 438512
rect 464396 438472 464402 438484
rect 508222 438472 508228 438484
rect 508280 438472 508286 438524
rect 382918 438404 382924 438456
rect 382976 438444 382982 438456
rect 402330 438444 402336 438456
rect 382976 438416 402336 438444
rect 382976 438404 382982 438416
rect 402330 438404 402336 438416
rect 402388 438404 402394 438456
rect 413278 438404 413284 438456
rect 413336 438444 413342 438456
rect 422938 438444 422944 438456
rect 413336 438416 422944 438444
rect 413336 438404 413342 438416
rect 422938 438404 422944 438416
rect 422996 438404 423002 438456
rect 460198 438404 460204 438456
rect 460256 438444 460262 438456
rect 503806 438444 503812 438456
rect 460256 438416 503812 438444
rect 460256 438404 460262 438416
rect 503806 438404 503812 438416
rect 503864 438404 503870 438456
rect 504358 438404 504364 438456
rect 504416 438444 504422 438456
rect 514110 438444 514116 438456
rect 504416 438416 514116 438444
rect 504416 438404 504422 438416
rect 514110 438404 514116 438416
rect 514168 438404 514174 438456
rect 388438 438336 388444 438388
rect 388496 438376 388502 438388
rect 415578 438376 415584 438388
rect 388496 438348 415584 438376
rect 388496 438336 388502 438348
rect 415578 438336 415584 438348
rect 415636 438336 415642 438388
rect 417418 438336 417424 438388
rect 417476 438376 417482 438388
rect 427354 438376 427360 438388
rect 417476 438348 427360 438376
rect 417476 438336 417482 438348
rect 427354 438336 427360 438348
rect 427412 438336 427418 438388
rect 446398 438336 446404 438388
rect 446456 438376 446462 438388
rect 494974 438376 494980 438388
rect 446456 438348 494980 438376
rect 446456 438336 446462 438348
rect 494974 438336 494980 438348
rect 495032 438336 495038 438388
rect 508498 438336 508504 438388
rect 508556 438376 508562 438388
rect 518526 438376 518532 438388
rect 508556 438348 518532 438376
rect 508556 438336 508562 438348
rect 518526 438336 518532 438348
rect 518584 438336 518590 438388
rect 358078 438268 358084 438320
rect 358136 438308 358142 438320
rect 419994 438308 420000 438320
rect 358136 438280 420000 438308
rect 358136 438268 358142 438280
rect 419994 438268 420000 438280
rect 420052 438268 420058 438320
rect 450538 438268 450544 438320
rect 450596 438308 450602 438320
rect 499574 438308 499580 438320
rect 450596 438280 499580 438308
rect 450596 438268 450602 438280
rect 499574 438268 499580 438280
rect 499632 438268 499638 438320
rect 501598 438268 501604 438320
rect 501656 438308 501662 438320
rect 509694 438308 509700 438320
rect 501656 438280 509700 438308
rect 501656 438268 501662 438280
rect 509694 438268 509700 438280
rect 509752 438268 509758 438320
rect 512638 438268 512644 438320
rect 512696 438308 512702 438320
rect 523034 438308 523040 438320
rect 512696 438280 523040 438308
rect 512696 438268 512702 438280
rect 523034 438268 523040 438280
rect 523092 438268 523098 438320
rect 392578 438200 392584 438252
rect 392636 438240 392642 438252
rect 469950 438240 469956 438252
rect 392636 438212 469956 438240
rect 392636 438200 392642 438212
rect 469950 438200 469956 438212
rect 470008 438200 470014 438252
rect 472618 438200 472624 438252
rect 472676 438240 472682 438252
rect 517054 438240 517060 438252
rect 472676 438212 517060 438240
rect 472676 438200 472682 438212
rect 517054 438200 517060 438212
rect 517112 438200 517118 438252
rect 518158 438200 518164 438252
rect 518216 438240 518222 438252
rect 527358 438240 527364 438252
rect 518216 438212 527364 438240
rect 518216 438200 518222 438212
rect 527358 438200 527364 438212
rect 527416 438200 527422 438252
rect 393958 438132 393964 438184
rect 394016 438172 394022 438184
rect 474366 438172 474372 438184
rect 394016 438144 474372 438172
rect 394016 438132 394022 438144
rect 474366 438132 474372 438144
rect 474424 438132 474430 438184
rect 475378 438132 475384 438184
rect 475436 438172 475442 438184
rect 521654 438172 521660 438184
rect 475436 438144 521660 438172
rect 475436 438132 475442 438144
rect 521654 438132 521660 438144
rect 521712 438132 521718 438184
rect 389818 437520 389824 437572
rect 389876 437560 389882 437572
rect 393498 437560 393504 437572
rect 389876 437532 393504 437560
rect 389876 437520 389882 437532
rect 393498 437520 393504 437532
rect 393556 437520 393562 437572
rect 497458 437520 497464 437572
rect 497516 437560 497522 437572
rect 500954 437560 500960 437572
rect 497516 437532 500960 437560
rect 497516 437520 497522 437532
rect 500954 437520 500960 437532
rect 501012 437520 501018 437572
rect 520918 437520 520924 437572
rect 520976 437560 520982 437572
rect 524414 437560 524420 437572
rect 520976 437532 524420 437560
rect 520976 437520 520982 437532
rect 524414 437520 524420 437532
rect 524472 437520 524478 437572
rect 389910 437452 389916 437504
rect 389968 437492 389974 437504
rect 390554 437492 390560 437504
rect 389968 437464 390560 437492
rect 389968 437452 389974 437464
rect 390554 437452 390560 437464
rect 390612 437452 390618 437504
rect 399478 437452 399484 437504
rect 399536 437492 399542 437504
rect 405274 437492 405280 437504
rect 399536 437464 405280 437492
rect 399536 437452 399542 437464
rect 405274 437452 405280 437464
rect 405332 437452 405338 437504
rect 443638 437452 443644 437504
rect 443696 437492 443702 437504
rect 445018 437492 445024 437504
rect 443696 437464 445024 437492
rect 443696 437452 443702 437464
rect 445018 437452 445024 437464
rect 445076 437452 445082 437504
rect 486418 437452 486424 437504
rect 486476 437492 486482 437504
rect 487614 437492 487620 437504
rect 486476 437464 487620 437492
rect 486476 437452 486482 437464
rect 487614 437452 487620 437464
rect 487672 437452 487678 437504
rect 490558 437452 490564 437504
rect 490616 437492 490622 437504
rect 492030 437492 492036 437504
rect 490616 437464 492036 437492
rect 490616 437452 490622 437464
rect 492030 437452 492036 437464
rect 492088 437452 492094 437504
rect 494698 437452 494704 437504
rect 494756 437492 494762 437504
rect 496446 437492 496452 437504
rect 494756 437464 496452 437492
rect 494756 437452 494762 437464
rect 496446 437452 496452 437464
rect 496504 437452 496510 437504
rect 500218 437452 500224 437504
rect 500276 437492 500282 437504
rect 505278 437492 505284 437504
rect 500276 437464 505284 437492
rect 500276 437452 500282 437464
rect 505278 437452 505284 437464
rect 505336 437452 505342 437504
rect 519538 437452 519544 437504
rect 519596 437492 519602 437504
rect 520274 437492 520280 437504
rect 519596 437464 520280 437492
rect 519596 437452 519602 437464
rect 520274 437452 520280 437464
rect 520332 437452 520338 437504
rect 522298 437452 522304 437504
rect 522356 437492 522362 437504
rect 528830 437492 528836 437504
rect 522356 437464 528836 437492
rect 522356 437452 522362 437464
rect 528830 437452 528836 437464
rect 528888 437452 528894 437504
rect 551278 431876 551284 431928
rect 551336 431916 551342 431928
rect 579798 431916 579804 431928
rect 551336 431888 579804 431916
rect 551336 431876 551342 431888
rect 579798 431876 579804 431888
rect 579856 431876 579862 431928
rect 558178 419432 558184 419484
rect 558236 419472 558242 419484
rect 580166 419472 580172 419484
rect 558236 419444 580172 419472
rect 558236 419432 558242 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 143442 396992 143448 397044
rect 143500 397032 143506 397044
rect 247034 397032 247040 397044
rect 143500 397004 247040 397032
rect 143500 396992 143506 397004
rect 247034 396992 247040 397004
rect 247092 396992 247098 397044
rect 142062 396924 142068 396976
rect 142120 396964 142126 396976
rect 245654 396964 245660 396976
rect 142120 396936 245660 396964
rect 142120 396924 142126 396936
rect 245654 396924 245660 396936
rect 245712 396924 245718 396976
rect 126882 396856 126888 396908
rect 126940 396896 126946 396908
rect 237374 396896 237380 396908
rect 126940 396868 237380 396896
rect 126940 396856 126946 396868
rect 237374 396856 237380 396868
rect 237432 396856 237438 396908
rect 124122 396788 124128 396840
rect 124180 396828 124186 396840
rect 235994 396828 236000 396840
rect 124180 396800 236000 396828
rect 124180 396788 124186 396800
rect 235994 396788 236000 396800
rect 236052 396788 236058 396840
rect 121362 396720 121368 396772
rect 121420 396760 121426 396772
rect 234614 396760 234620 396772
rect 121420 396732 234620 396760
rect 121420 396720 121426 396732
rect 234614 396720 234620 396732
rect 234672 396720 234678 396772
rect 118602 395632 118608 395684
rect 118660 395672 118666 395684
rect 233234 395672 233240 395684
rect 118660 395644 233240 395672
rect 118660 395632 118666 395644
rect 233234 395632 233240 395644
rect 233292 395632 233298 395684
rect 117222 395564 117228 395616
rect 117280 395604 117286 395616
rect 231854 395604 231860 395616
rect 117280 395576 231860 395604
rect 117280 395564 117286 395576
rect 231854 395564 231860 395576
rect 231912 395564 231918 395616
rect 114462 395496 114468 395548
rect 114520 395536 114526 395548
rect 230474 395536 230480 395548
rect 114520 395508 230480 395536
rect 114520 395496 114526 395508
rect 230474 395496 230480 395508
rect 230532 395496 230538 395548
rect 111702 395428 111708 395480
rect 111760 395468 111766 395480
rect 229094 395468 229100 395480
rect 111760 395440 229100 395468
rect 111760 395428 111766 395440
rect 229094 395428 229100 395440
rect 229152 395428 229158 395480
rect 108942 395360 108948 395412
rect 109000 395400 109006 395412
rect 227714 395400 227720 395412
rect 109000 395372 227720 395400
rect 109000 395360 109006 395372
rect 227714 395360 227720 395372
rect 227772 395360 227778 395412
rect 106182 395292 106188 395344
rect 106240 395332 106246 395344
rect 226334 395332 226340 395344
rect 106240 395304 226340 395332
rect 106240 395292 106246 395304
rect 226334 395292 226340 395304
rect 226392 395292 226398 395344
rect 157334 394272 157340 394324
rect 157392 394312 157398 394324
rect 270494 394312 270500 394324
rect 157392 394284 270500 394312
rect 157392 394272 157398 394284
rect 270494 394272 270500 394284
rect 270552 394272 270558 394324
rect 104802 394204 104808 394256
rect 104860 394244 104866 394256
rect 223574 394244 223580 394256
rect 104860 394216 223580 394244
rect 104860 394204 104866 394216
rect 223574 394204 223580 394216
rect 223632 394204 223638 394256
rect 102042 394136 102048 394188
rect 102100 394176 102106 394188
rect 222194 394176 222200 394188
rect 102100 394148 222200 394176
rect 102100 394136 102106 394148
rect 222194 394136 222200 394148
rect 222252 394136 222258 394188
rect 99282 394068 99288 394120
rect 99340 394108 99346 394120
rect 220814 394108 220820 394120
rect 99340 394080 220820 394108
rect 99340 394068 99346 394080
rect 220814 394068 220820 394080
rect 220872 394068 220878 394120
rect 96522 394000 96528 394052
rect 96580 394040 96586 394052
rect 219434 394040 219440 394052
rect 96580 394012 219440 394040
rect 96580 394000 96586 394012
rect 219434 394000 219440 394012
rect 219492 394000 219498 394052
rect 93762 393932 93768 393984
rect 93820 393972 93826 393984
rect 218054 393972 218060 393984
rect 93820 393944 218060 393972
rect 93820 393932 93826 393944
rect 218054 393932 218060 393944
rect 218112 393932 218118 393984
rect 149054 392980 149060 393032
rect 149112 393020 149118 393032
rect 255314 393020 255320 393032
rect 149112 392992 255320 393020
rect 149112 392980 149118 392992
rect 255314 392980 255320 392992
rect 255372 392980 255378 393032
rect 150434 392912 150440 392964
rect 150492 392952 150498 392964
rect 258258 392952 258264 392964
rect 150492 392924 258264 392952
rect 150492 392912 150498 392924
rect 258258 392912 258264 392924
rect 258316 392912 258322 392964
rect 151814 392844 151820 392896
rect 151872 392884 151878 392896
rect 260834 392884 260840 392896
rect 151872 392856 260840 392884
rect 151872 392844 151878 392856
rect 260834 392844 260840 392856
rect 260892 392844 260898 392896
rect 153194 392776 153200 392828
rect 153252 392816 153258 392828
rect 263594 392816 263600 392828
rect 153252 392788 263600 392816
rect 153252 392776 153258 392788
rect 263594 392776 263600 392788
rect 263652 392776 263658 392828
rect 154574 392708 154580 392760
rect 154632 392748 154638 392760
rect 264974 392748 264980 392760
rect 154632 392720 264980 392748
rect 154632 392708 154638 392720
rect 264974 392708 264980 392720
rect 265032 392708 265038 392760
rect 155954 392640 155960 392692
rect 156012 392680 156018 392692
rect 268102 392680 268108 392692
rect 156012 392652 268108 392680
rect 156012 392640 156018 392652
rect 268102 392640 268108 392652
rect 268160 392640 268166 392692
rect 71314 392572 71320 392624
rect 71372 392612 71378 392624
rect 205634 392612 205640 392624
rect 71372 392584 205640 392612
rect 71372 392572 71378 392584
rect 205634 392572 205640 392584
rect 205692 392572 205698 392624
rect 147674 391620 147680 391672
rect 147732 391660 147738 391672
rect 252554 391660 252560 391672
rect 147732 391632 252560 391660
rect 147732 391620 147738 391632
rect 252554 391620 252560 391632
rect 252612 391620 252618 391672
rect 158714 391552 158720 391604
rect 158772 391592 158778 391604
rect 273254 391592 273260 391604
rect 158772 391564 273260 391592
rect 158772 391552 158778 391564
rect 273254 391552 273260 391564
rect 273312 391552 273318 391604
rect 161474 391484 161480 391536
rect 161532 391524 161538 391536
rect 277946 391524 277952 391536
rect 161532 391496 277952 391524
rect 161532 391484 161538 391496
rect 277946 391484 277952 391496
rect 278004 391484 278010 391536
rect 160094 391416 160100 391468
rect 160152 391456 160158 391468
rect 276014 391456 276020 391468
rect 160152 391428 276020 391456
rect 160152 391416 160158 391428
rect 276014 391416 276020 391428
rect 276072 391416 276078 391468
rect 162854 391348 162860 391400
rect 162912 391388 162918 391400
rect 280154 391388 280160 391400
rect 162912 391360 280160 391388
rect 162912 391348 162918 391360
rect 280154 391348 280160 391360
rect 280212 391348 280218 391400
rect 68738 391280 68744 391332
rect 68796 391320 68802 391332
rect 204254 391320 204260 391332
rect 68796 391292 204260 391320
rect 68796 391280 68802 391292
rect 204254 391280 204260 391292
rect 204312 391280 204318 391332
rect 189074 391212 189080 391264
rect 189132 391252 189138 391264
rect 325878 391252 325884 391264
rect 189132 391224 325884 391252
rect 189132 391212 189138 391224
rect 325878 391212 325884 391224
rect 325936 391212 325942 391264
rect 159818 390192 159824 390244
rect 159876 390232 159882 390244
rect 191834 390232 191840 390244
rect 159876 390204 191840 390232
rect 159876 390192 159882 390204
rect 191834 390192 191840 390204
rect 191892 390192 191898 390244
rect 158530 390124 158536 390176
rect 158588 390164 158594 390176
rect 193214 390164 193220 390176
rect 158588 390136 193220 390164
rect 158588 390124 158594 390136
rect 193214 390124 193220 390136
rect 193272 390124 193278 390176
rect 144914 390056 144920 390108
rect 144972 390096 144978 390108
rect 248506 390096 248512 390108
rect 144972 390068 248512 390096
rect 144972 390056 144978 390068
rect 248506 390056 248512 390068
rect 248564 390056 248570 390108
rect 186314 389988 186320 390040
rect 186372 390028 186378 390040
rect 320174 390028 320180 390040
rect 186372 390000 320180 390028
rect 186372 389988 186378 390000
rect 320174 389988 320180 390000
rect 320232 389988 320238 390040
rect 132494 389920 132500 389972
rect 132552 389960 132558 389972
rect 338114 389960 338120 389972
rect 132552 389932 338120 389960
rect 132552 389920 132558 389932
rect 338114 389920 338120 389932
rect 338172 389920 338178 389972
rect 131114 389852 131120 389904
rect 131172 389892 131178 389904
rect 339494 389892 339500 389904
rect 131172 389864 339500 389892
rect 131172 389852 131178 389864
rect 339494 389852 339500 389864
rect 339552 389852 339558 389904
rect 129734 389784 129740 389836
rect 129792 389824 129798 389836
rect 359274 389824 359280 389836
rect 129792 389796 359280 389824
rect 129792 389784 129798 389796
rect 359274 389784 359280 389796
rect 359332 389784 359338 389836
rect 176654 388832 176660 388884
rect 176712 388872 176718 388884
rect 304994 388872 305000 388884
rect 176712 388844 305000 388872
rect 176712 388832 176718 388844
rect 304994 388832 305000 388844
rect 305052 388832 305058 388884
rect 178034 388764 178040 388816
rect 178092 388804 178098 388816
rect 307754 388804 307760 388816
rect 178092 388776 307760 388804
rect 178092 388764 178098 388776
rect 307754 388764 307760 388776
rect 307812 388764 307818 388816
rect 179414 388696 179420 388748
rect 179472 388736 179478 388748
rect 310514 388736 310520 388748
rect 179472 388708 310520 388736
rect 179472 388696 179478 388708
rect 310514 388696 310520 388708
rect 310572 388696 310578 388748
rect 180794 388628 180800 388680
rect 180852 388668 180858 388680
rect 313274 388668 313280 388680
rect 180852 388640 313280 388668
rect 180852 388628 180858 388640
rect 313274 388628 313280 388640
rect 313332 388628 313338 388680
rect 183554 388560 183560 388612
rect 183612 388600 183618 388612
rect 317414 388600 317420 388612
rect 183612 388572 317420 388600
rect 183612 388560 183618 388572
rect 317414 388560 317420 388572
rect 317472 388560 317478 388612
rect 182174 388492 182180 388544
rect 182232 388532 182238 388544
rect 316034 388532 316040 388544
rect 182232 388504 316040 388532
rect 182232 388492 182238 388504
rect 316034 388492 316040 388504
rect 316092 388492 316098 388544
rect 187694 388424 187700 388476
rect 187752 388464 187758 388476
rect 322934 388464 322940 388476
rect 187752 388436 322940 388464
rect 187752 388424 187758 388436
rect 322934 388424 322940 388436
rect 322992 388424 322998 388476
rect 146294 387676 146300 387728
rect 146352 387716 146358 387728
rect 249794 387716 249800 387728
rect 146352 387688 249800 387716
rect 146352 387676 146358 387688
rect 249794 387676 249800 387688
rect 249852 387676 249858 387728
rect 164234 387608 164240 387660
rect 164292 387648 164298 387660
rect 282914 387648 282920 387660
rect 164292 387620 282920 387648
rect 164292 387608 164298 387620
rect 282914 387608 282920 387620
rect 282972 387608 282978 387660
rect 165614 387540 165620 387592
rect 165672 387580 165678 387592
rect 285674 387580 285680 387592
rect 165672 387552 285680 387580
rect 165672 387540 165678 387552
rect 285674 387540 285680 387552
rect 285732 387540 285738 387592
rect 166994 387472 167000 387524
rect 167052 387512 167058 387524
rect 288434 387512 288440 387524
rect 167052 387484 288440 387512
rect 167052 387472 167058 387484
rect 288434 387472 288440 387484
rect 288492 387472 288498 387524
rect 168374 387404 168380 387456
rect 168432 387444 168438 387456
rect 289814 387444 289820 387456
rect 168432 387416 289820 387444
rect 168432 387404 168438 387416
rect 289814 387404 289820 387416
rect 289872 387404 289878 387456
rect 169754 387336 169760 387388
rect 169812 387376 169818 387388
rect 292574 387376 292580 387388
rect 169812 387348 292580 387376
rect 169812 387336 169818 387348
rect 292574 387336 292580 387348
rect 292632 387336 292638 387388
rect 171134 387268 171140 387320
rect 171192 387308 171198 387320
rect 295334 387308 295340 387320
rect 171192 387280 295340 387308
rect 171192 387268 171198 387280
rect 295334 387268 295340 387280
rect 295392 387268 295398 387320
rect 172514 387200 172520 387252
rect 172572 387240 172578 387252
rect 298094 387240 298100 387252
rect 172572 387212 298100 387240
rect 172572 387200 172578 387212
rect 298094 387200 298100 387212
rect 298152 387200 298158 387252
rect 175274 387132 175280 387184
rect 175332 387172 175338 387184
rect 302234 387172 302240 387184
rect 175332 387144 302240 387172
rect 175332 387132 175338 387144
rect 302234 387132 302240 387144
rect 302292 387132 302298 387184
rect 173894 387064 173900 387116
rect 173952 387104 173958 387116
rect 300854 387104 300860 387116
rect 173952 387076 300860 387104
rect 173952 387064 173958 387076
rect 300854 387064 300860 387076
rect 300912 387064 300918 387116
rect 78490 386316 78496 386368
rect 78548 386356 78554 386368
rect 80698 386356 80704 386368
rect 78548 386328 80704 386356
rect 78548 386316 78554 386328
rect 80698 386316 80704 386328
rect 80756 386316 80762 386368
rect 89162 386316 89168 386368
rect 89220 386356 89226 386368
rect 90358 386356 90364 386368
rect 89220 386328 90364 386356
rect 89220 386316 89226 386328
rect 90358 386316 90364 386328
rect 90416 386316 90422 386368
rect 133690 386316 133696 386368
rect 133748 386356 133754 386368
rect 134518 386356 134524 386368
rect 133748 386328 134524 386356
rect 133748 386316 133754 386328
rect 134518 386316 134524 386328
rect 134576 386316 134582 386368
rect 138474 386316 138480 386368
rect 138532 386356 138538 386368
rect 140038 386356 140044 386368
rect 138532 386328 140044 386356
rect 138532 386316 138538 386328
rect 140038 386316 140044 386328
rect 140096 386316 140102 386368
rect 146202 386316 146208 386368
rect 146260 386356 146266 386368
rect 155218 386356 155224 386368
rect 146260 386328 155224 386356
rect 146260 386316 146266 386328
rect 155218 386316 155224 386328
rect 155276 386316 155282 386368
rect 73890 386248 73896 386300
rect 73948 386288 73954 386300
rect 79318 386288 79324 386300
rect 73948 386260 79324 386288
rect 73948 386248 73954 386260
rect 79318 386248 79324 386260
rect 79376 386248 79382 386300
rect 81066 386248 81072 386300
rect 81124 386288 81130 386300
rect 211154 386288 211160 386300
rect 81124 386260 211160 386288
rect 81124 386248 81130 386260
rect 211154 386248 211160 386260
rect 211212 386248 211218 386300
rect 86494 386180 86500 386232
rect 86552 386220 86558 386232
rect 213914 386220 213920 386232
rect 86552 386192 213920 386220
rect 86552 386180 86558 386192
rect 213914 386180 213920 386192
rect 213972 386180 213978 386232
rect 92106 386112 92112 386164
rect 92164 386152 92170 386164
rect 216674 386152 216680 386164
rect 92164 386124 216680 386152
rect 92164 386112 92170 386124
rect 216674 386112 216680 386124
rect 216732 386112 216738 386164
rect 131022 386044 131028 386096
rect 131080 386084 131086 386096
rect 218882 386084 218888 386096
rect 131080 386056 218888 386084
rect 131080 386044 131086 386056
rect 218882 386044 218888 386056
rect 218940 386044 218946 386096
rect 136082 385976 136088 386028
rect 136140 386016 136146 386028
rect 220078 386016 220084 386028
rect 136140 385988 220084 386016
rect 136140 385976 136146 385988
rect 220078 385976 220084 385988
rect 220136 385976 220142 386028
rect 128630 385908 128636 385960
rect 128688 385948 128694 385960
rect 152458 385948 152464 385960
rect 128688 385920 152464 385948
rect 128688 385908 128694 385920
rect 152458 385908 152464 385920
rect 152516 385908 152522 385960
rect 77202 385840 77208 385892
rect 77260 385880 77266 385892
rect 208394 385880 208400 385892
rect 77260 385852 208400 385880
rect 77260 385840 77266 385852
rect 208394 385840 208400 385852
rect 208452 385840 208458 385892
rect 350994 385636 351000 385688
rect 351052 385676 351058 385688
rect 380894 385676 380900 385688
rect 351052 385648 380900 385676
rect 351052 385636 351058 385648
rect 380894 385636 380900 385648
rect 380952 385636 380958 385688
rect 83642 385092 83648 385144
rect 83700 385132 83706 385144
rect 86218 385132 86224 385144
rect 83700 385104 86224 385132
rect 83700 385092 83706 385104
rect 86218 385092 86224 385104
rect 86276 385092 86282 385144
rect 170858 384616 170864 384668
rect 170916 384656 170922 384668
rect 177298 384656 177304 384668
rect 170916 384628 177304 384656
rect 170916 384616 170922 384628
rect 177298 384616 177304 384628
rect 177356 384616 177362 384668
rect 217870 384616 217876 384668
rect 217928 384656 217934 384668
rect 350994 384656 351000 384668
rect 217928 384628 351000 384656
rect 217928 384616 217934 384628
rect 350994 384616 351000 384628
rect 351052 384616 351058 384668
rect 139394 384548 139400 384600
rect 139452 384588 139458 384600
rect 358814 384588 358820 384600
rect 139452 384560 358820 384588
rect 139452 384548 139458 384560
rect 358814 384548 358820 384560
rect 358872 384548 358878 384600
rect 138014 384480 138020 384532
rect 138072 384520 138078 384532
rect 358906 384520 358912 384532
rect 138072 384492 358912 384520
rect 138072 384480 138078 384492
rect 358906 384480 358912 384492
rect 358964 384480 358970 384532
rect 136634 384412 136640 384464
rect 136692 384452 136698 384464
rect 358998 384452 359004 384464
rect 136692 384424 359004 384452
rect 136692 384412 136698 384424
rect 358998 384412 359004 384424
rect 359056 384412 359062 384464
rect 135254 384344 135260 384396
rect 135312 384384 135318 384396
rect 359090 384384 359096 384396
rect 135312 384356 359096 384384
rect 135312 384344 135318 384356
rect 359090 384344 359096 384356
rect 359148 384344 359154 384396
rect 133874 384276 133880 384328
rect 133932 384316 133938 384328
rect 359182 384316 359188 384328
rect 133932 384288 359188 384316
rect 133932 384276 133938 384288
rect 359182 384276 359188 384288
rect 359240 384276 359246 384328
rect 178678 379448 178684 379500
rect 178736 379488 178742 379500
rect 190454 379488 190460 379500
rect 178736 379460 190460 379488
rect 178736 379448 178742 379460
rect 190454 379448 190460 379460
rect 190512 379448 190518 379500
rect 548518 379448 548524 379500
rect 548576 379488 548582 379500
rect 580166 379488 580172 379500
rect 548576 379460 580172 379488
rect 548576 379448 548582 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 556798 365644 556804 365696
rect 556856 365684 556862 365696
rect 580166 365684 580172 365696
rect 556856 365656 580172 365684
rect 556856 365644 556862 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 176654 336744 176660 336796
rect 176712 336784 176718 336796
rect 216674 336784 216680 336796
rect 176712 336756 216680 336784
rect 176712 336744 176718 336756
rect 216674 336744 216680 336756
rect 216732 336744 216738 336796
rect 178678 320084 178684 320136
rect 178736 320124 178742 320136
rect 194594 320124 194600 320136
rect 178736 320096 194600 320124
rect 178736 320084 178742 320096
rect 194594 320084 194600 320096
rect 194652 320084 194658 320136
rect 178954 318724 178960 318776
rect 179012 318764 179018 318776
rect 195974 318764 195980 318776
rect 179012 318736 195980 318764
rect 179012 318724 179018 318736
rect 195974 318724 195980 318736
rect 196032 318724 196038 318776
rect 178954 317364 178960 317416
rect 179012 317404 179018 317416
rect 197354 317404 197360 317416
rect 179012 317376 197360 317404
rect 179012 317364 179018 317376
rect 197354 317364 197360 317376
rect 197412 317364 197418 317416
rect 178586 315936 178592 315988
rect 178644 315976 178650 315988
rect 198734 315976 198740 315988
rect 178644 315948 198740 315976
rect 178644 315936 178650 315948
rect 198734 315936 198740 315948
rect 198792 315936 198798 315988
rect 178678 314576 178684 314628
rect 178736 314616 178742 314628
rect 200114 314616 200120 314628
rect 178736 314588 200120 314616
rect 178736 314576 178742 314588
rect 200114 314576 200120 314588
rect 200172 314576 200178 314628
rect 182818 309136 182824 309188
rect 182876 309176 182882 309188
rect 216674 309176 216680 309188
rect 182876 309148 216680 309176
rect 182876 309136 182882 309148
rect 216674 309136 216680 309148
rect 216732 309136 216738 309188
rect 177298 309068 177304 309120
rect 177356 309108 177362 309120
rect 216766 309108 216772 309120
rect 177356 309080 216772 309108
rect 177356 309068 177362 309080
rect 216766 309068 216772 309080
rect 216824 309068 216830 309120
rect 39114 299412 39120 299464
rect 39172 299452 39178 299464
rect 39942 299452 39948 299464
rect 39172 299424 39948 299452
rect 39172 299412 39178 299424
rect 39942 299412 39948 299424
rect 40000 299452 40006 299464
rect 177298 299452 177304 299464
rect 40000 299424 177304 299452
rect 40000 299412 40006 299424
rect 177298 299412 177304 299424
rect 177356 299412 177362 299464
rect 163222 298868 163228 298920
rect 163280 298908 163286 298920
rect 201494 298908 201500 298920
rect 163280 298880 201500 298908
rect 163280 298868 163286 298880
rect 201494 298868 201500 298880
rect 201552 298868 201558 298920
rect 163406 298732 163412 298784
rect 163464 298772 163470 298784
rect 202874 298772 202880 298784
rect 163464 298744 202880 298772
rect 163464 298732 163470 298744
rect 202874 298732 202880 298744
rect 202932 298732 202938 298784
rect 218698 298052 218704 298104
rect 218756 298092 218762 298104
rect 343358 298092 343364 298104
rect 218756 298064 343364 298092
rect 218756 298052 218762 298064
rect 343358 298052 343364 298064
rect 343416 298052 343422 298104
rect 136082 297984 136088 298036
rect 136140 298024 136146 298036
rect 140038 298024 140044 298036
rect 136140 297996 140044 298024
rect 136140 297984 136146 297996
rect 140038 297984 140044 297996
rect 140096 297984 140102 298036
rect 218790 297984 218796 298036
rect 218848 298024 218854 298036
rect 343174 298024 343180 298036
rect 218848 297996 343180 298024
rect 218848 297984 218854 297996
rect 343174 297984 343180 297996
rect 343232 297984 343238 298036
rect 264330 297916 264336 297968
rect 264388 297956 264394 297968
rect 265342 297956 265348 297968
rect 264388 297928 265348 297956
rect 264388 297916 264394 297928
rect 265342 297916 265348 297928
rect 265400 297916 265406 297968
rect 275278 297916 275284 297968
rect 275336 297956 275342 297968
rect 276750 297956 276756 297968
rect 275336 297928 276756 297956
rect 275336 297916 275342 297928
rect 276750 297916 276756 297928
rect 276808 297916 276814 297968
rect 282178 297916 282184 297968
rect 282236 297956 282242 297968
rect 285950 297956 285956 297968
rect 282236 297928 285956 297956
rect 282236 297916 282242 297928
rect 285950 297916 285956 297928
rect 286008 297916 286014 297968
rect 287698 297916 287704 297968
rect 287756 297956 287762 297968
rect 295334 297956 295340 297968
rect 287756 297928 295340 297956
rect 287756 297916 287762 297928
rect 295334 297916 295340 297928
rect 295392 297916 295398 297968
rect 68830 297848 68836 297900
rect 68888 297888 68894 297900
rect 69658 297888 69664 297900
rect 68888 297860 69664 297888
rect 68888 297848 68894 297860
rect 69658 297848 69664 297860
rect 69716 297848 69722 297900
rect 77202 297304 77208 297356
rect 77260 297344 77266 297356
rect 259546 297344 259552 297356
rect 77260 297316 259552 297344
rect 77260 297304 77266 297316
rect 259546 297304 259552 297316
rect 259604 297304 259610 297356
rect 203518 297236 203524 297288
rect 203576 297276 203582 297288
rect 238110 297276 238116 297288
rect 203576 297248 238116 297276
rect 203576 297236 203582 297248
rect 238110 297236 238116 297248
rect 238168 297236 238174 297288
rect 108574 297168 108580 297220
rect 108632 297208 108638 297220
rect 125870 297208 125876 297220
rect 108632 297180 125876 297208
rect 108632 297168 108638 297180
rect 125870 297168 125876 297180
rect 125928 297168 125934 297220
rect 141050 297168 141056 297220
rect 141108 297208 141114 297220
rect 162118 297208 162124 297220
rect 141108 297180 162124 297208
rect 141108 297168 141114 297180
rect 162118 297168 162124 297180
rect 162176 297168 162182 297220
rect 202138 297168 202144 297220
rect 202196 297208 202202 297220
rect 276014 297208 276020 297220
rect 202196 297180 276020 297208
rect 202196 297168 202202 297180
rect 276014 297168 276020 297180
rect 276072 297168 276078 297220
rect 108942 297100 108948 297152
rect 109000 297140 109006 297152
rect 251542 297140 251548 297152
rect 109000 297112 251548 297140
rect 109000 297100 109006 297112
rect 251542 297100 251548 297112
rect 251600 297100 251606 297152
rect 108850 297032 108856 297084
rect 108908 297072 108914 297084
rect 259454 297072 259460 297084
rect 108908 297044 259460 297072
rect 108908 297032 108914 297044
rect 259454 297032 259460 297044
rect 259512 297032 259518 297084
rect 302878 297032 302884 297084
rect 302936 297072 302942 297084
rect 315758 297072 315764 297084
rect 302936 297044 315764 297072
rect 302936 297032 302942 297044
rect 315758 297032 315764 297044
rect 315816 297032 315822 297084
rect 108666 296964 108672 297016
rect 108724 297004 108730 297016
rect 269758 297004 269764 297016
rect 108724 296976 269764 297004
rect 108724 296964 108730 296976
rect 269758 296964 269764 296976
rect 269816 296964 269822 297016
rect 294598 296964 294604 297016
rect 294656 297004 294662 297016
rect 302326 297004 302332 297016
rect 294656 296976 302332 297004
rect 294656 296964 294662 296976
rect 302326 296964 302332 296976
rect 302384 296964 302390 297016
rect 305638 296964 305644 297016
rect 305696 297004 305702 297016
rect 320910 297004 320916 297016
rect 305696 296976 320916 297004
rect 305696 296964 305702 296976
rect 320910 296964 320916 296976
rect 320968 296964 320974 297016
rect 86218 296896 86224 296948
rect 86276 296936 86282 296948
rect 259454 296936 259460 296948
rect 86276 296908 259460 296936
rect 86276 296896 86282 296908
rect 259454 296896 259460 296908
rect 259512 296896 259518 296948
rect 289078 296896 289084 296948
rect 289136 296936 289142 296948
rect 298462 296936 298468 296948
rect 289136 296908 298468 296936
rect 289136 296896 289142 296908
rect 298462 296896 298468 296908
rect 298520 296896 298526 296948
rect 300118 296896 300124 296948
rect 300176 296936 300182 296948
rect 310974 296936 310980 296948
rect 300176 296908 310980 296936
rect 300176 296896 300182 296908
rect 310974 296896 310980 296908
rect 311032 296896 311038 296948
rect 83366 296828 83372 296880
rect 83424 296868 83430 296880
rect 259730 296868 259736 296880
rect 83424 296840 259736 296868
rect 83424 296828 83430 296840
rect 259730 296828 259736 296840
rect 259788 296828 259794 296880
rect 295978 296828 295984 296880
rect 296036 296868 296042 296880
rect 305086 296868 305092 296880
rect 296036 296840 305092 296868
rect 296036 296828 296042 296840
rect 305086 296828 305092 296840
rect 305144 296828 305150 296880
rect 80698 296760 80704 296812
rect 80756 296800 80762 296812
rect 259638 296800 259644 296812
rect 80756 296772 259644 296800
rect 80756 296760 80762 296772
rect 259638 296760 259644 296772
rect 259696 296760 259702 296812
rect 286318 296760 286324 296812
rect 286376 296800 286382 296812
rect 289998 296800 290004 296812
rect 286376 296772 290004 296800
rect 286376 296760 286382 296772
rect 289998 296760 290004 296772
rect 290056 296760 290062 296812
rect 291838 296760 291844 296812
rect 291896 296800 291902 296812
rect 300854 296800 300860 296812
rect 291896 296772 300860 296800
rect 291896 296760 291902 296772
rect 300854 296760 300860 296772
rect 300912 296760 300918 296812
rect 304258 296760 304264 296812
rect 304316 296800 304322 296812
rect 317414 296800 317420 296812
rect 304316 296772 317420 296800
rect 304316 296760 304322 296772
rect 317414 296760 317420 296772
rect 317472 296760 317478 296812
rect 108758 296692 108764 296744
rect 108816 296732 108822 296744
rect 117406 296732 117412 296744
rect 108816 296704 117412 296732
rect 108816 296692 108822 296704
rect 117406 296692 117412 296704
rect 117464 296692 117470 296744
rect 129642 296692 129648 296744
rect 129700 296732 129706 296744
rect 137278 296732 137284 296744
rect 129700 296704 137284 296732
rect 129700 296692 129706 296704
rect 137278 296692 137284 296704
rect 137336 296692 137342 296744
rect 264238 296692 264244 296744
rect 264296 296732 264302 296744
rect 268010 296732 268016 296744
rect 264296 296704 268016 296732
rect 264296 296692 264302 296704
rect 268010 296692 268016 296704
rect 268068 296692 268074 296744
rect 284938 296692 284944 296744
rect 284996 296732 285002 296744
rect 287606 296732 287612 296744
rect 284996 296704 287612 296732
rect 284996 296692 285002 296704
rect 287606 296692 287612 296704
rect 287664 296692 287670 296744
rect 298738 296692 298744 296744
rect 298796 296732 298802 296744
rect 308582 296732 308588 296744
rect 298796 296704 308588 296732
rect 298796 296692 298802 296704
rect 308582 296692 308588 296704
rect 308640 296692 308646 296744
rect 205634 296012 205640 296064
rect 205692 296052 205698 296064
rect 261110 296052 261116 296064
rect 205692 296024 261116 296052
rect 205692 296012 205698 296024
rect 261110 296012 261116 296024
rect 261168 296012 261174 296064
rect 198734 295944 198740 295996
rect 198792 295984 198798 295996
rect 260190 295984 260196 295996
rect 198792 295956 260196 295984
rect 198792 295944 198798 295956
rect 260190 295944 260196 295956
rect 260248 295944 260254 295996
rect 160094 242156 160100 242208
rect 160152 242196 160158 242208
rect 260926 242196 260932 242208
rect 160152 242168 260932 242196
rect 160152 242156 160158 242168
rect 260926 242156 260932 242168
rect 260984 242156 260990 242208
rect 191834 240932 191840 240984
rect 191892 240972 191898 240984
rect 280154 240972 280160 240984
rect 191892 240944 280160 240972
rect 191892 240932 191898 240944
rect 280154 240932 280160 240944
rect 280212 240932 280218 240984
rect 109218 240864 109224 240916
rect 109276 240904 109282 240916
rect 292574 240904 292580 240916
rect 109276 240876 292580 240904
rect 109276 240864 109282 240876
rect 292574 240864 292580 240876
rect 292632 240864 292638 240916
rect 73062 240796 73068 240848
rect 73120 240836 73126 240848
rect 260190 240836 260196 240848
rect 73120 240808 260196 240836
rect 73120 240796 73126 240808
rect 260190 240796 260196 240808
rect 260248 240796 260254 240848
rect 109586 240728 109592 240780
rect 109644 240768 109650 240780
rect 313274 240768 313280 240780
rect 109644 240740 313280 240768
rect 109644 240728 109650 240740
rect 313274 240728 313280 240740
rect 313332 240728 313338 240780
rect 71682 239368 71688 239420
rect 71740 239408 71746 239420
rect 260098 239408 260104 239420
rect 71740 239380 260104 239408
rect 71740 239368 71746 239380
rect 260098 239368 260104 239380
rect 260156 239368 260162 239420
rect 89622 238076 89628 238128
rect 89680 238116 89686 238128
rect 229830 238116 229836 238128
rect 89680 238088 229836 238116
rect 89680 238076 89686 238088
rect 229830 238076 229836 238088
rect 229888 238076 229894 238128
rect 90910 238008 90916 238060
rect 90968 238048 90974 238060
rect 233326 238048 233332 238060
rect 90968 238020 233332 238048
rect 90968 238008 90974 238020
rect 233326 238008 233332 238020
rect 233384 238008 233390 238060
rect 174722 236988 174728 237040
rect 174780 237028 174786 237040
rect 251358 237028 251364 237040
rect 174780 237000 251364 237028
rect 174780 236988 174786 237000
rect 251358 236988 251364 237000
rect 251416 236988 251422 237040
rect 167730 236920 167736 236972
rect 167788 236960 167794 236972
rect 249794 236960 249800 236972
rect 167788 236932 249800 236960
rect 167788 236920 167794 236932
rect 249794 236920 249800 236932
rect 249852 236920 249858 236972
rect 157242 236852 157248 236904
rect 157300 236892 157306 236904
rect 248414 236892 248420 236904
rect 157300 236864 248420 236892
rect 157300 236852 157306 236864
rect 248414 236852 248420 236864
rect 248472 236852 248478 236904
rect 82722 236784 82728 236836
rect 82780 236824 82786 236836
rect 208946 236824 208952 236836
rect 82780 236796 208952 236824
rect 82780 236784 82786 236796
rect 208946 236784 208952 236796
rect 209004 236784 209010 236836
rect 244182 236784 244188 236836
rect 244240 236824 244246 236836
rect 273438 236824 273444 236836
rect 244240 236796 273444 236824
rect 244240 236784 244246 236796
rect 273438 236784 273444 236796
rect 273496 236784 273502 236836
rect 84010 236716 84016 236768
rect 84068 236756 84074 236768
rect 222930 236756 222936 236768
rect 84068 236728 222936 236756
rect 84068 236716 84074 236728
rect 222930 236716 222936 236728
rect 222988 236716 222994 236768
rect 240962 236716 240968 236768
rect 241020 236756 241026 236768
rect 271874 236756 271880 236768
rect 241020 236728 271880 236756
rect 241020 236716 241026 236728
rect 271874 236716 271880 236728
rect 271932 236716 271938 236768
rect 77110 236648 77116 236700
rect 77168 236688 77174 236700
rect 260282 236688 260288 236700
rect 77168 236660 260288 236688
rect 77168 236648 77174 236660
rect 260282 236648 260288 236660
rect 260340 236648 260346 236700
rect 38930 235560 38936 235612
rect 38988 235600 38994 235612
rect 111334 235600 111340 235612
rect 38988 235572 111340 235600
rect 38988 235560 38994 235572
rect 111334 235560 111340 235572
rect 111392 235560 111398 235612
rect 188614 235560 188620 235612
rect 188672 235600 188678 235612
rect 258166 235600 258172 235612
rect 188672 235572 258172 235600
rect 188672 235560 188678 235572
rect 258166 235560 258172 235572
rect 258224 235560 258230 235612
rect 79962 235492 79968 235544
rect 80020 235532 80026 235544
rect 194962 235532 194968 235544
rect 80020 235504 194968 235532
rect 80020 235492 80026 235504
rect 194962 235492 194968 235504
rect 195020 235492 195026 235544
rect 216582 235492 216588 235544
rect 216640 235532 216646 235544
rect 262214 235532 262220 235544
rect 216640 235504 262220 235532
rect 216640 235492 216646 235504
rect 262214 235492 262220 235504
rect 262272 235492 262278 235544
rect 109034 235424 109040 235476
rect 109092 235464 109098 235476
rect 255314 235464 255320 235476
rect 109092 235436 255320 235464
rect 109092 235424 109098 235436
rect 255314 235424 255320 235436
rect 255372 235424 255378 235476
rect 109126 235356 109132 235408
rect 109184 235396 109190 235408
rect 256694 235396 256700 235408
rect 109184 235368 256700 235396
rect 109184 235356 109190 235368
rect 256694 235356 256700 235368
rect 256752 235356 256758 235408
rect 109310 235288 109316 235340
rect 109368 235328 109374 235340
rect 265066 235328 265072 235340
rect 109368 235300 265072 235328
rect 109368 235288 109374 235300
rect 265066 235288 265072 235300
rect 265124 235288 265130 235340
rect 109402 235220 109408 235272
rect 109460 235260 109466 235272
rect 267826 235260 267832 235272
rect 109460 235232 267832 235260
rect 109460 235220 109466 235232
rect 267826 235220 267832 235232
rect 267884 235220 267890 235272
rect 57882 234132 57888 234184
rect 57940 234172 57946 234184
rect 132586 234172 132592 234184
rect 57940 234144 132592 234172
rect 57940 234132 57946 234144
rect 132586 234132 132592 234144
rect 132644 234132 132650 234184
rect 136358 234132 136364 234184
rect 136416 234172 136422 234184
rect 217502 234172 217508 234184
rect 136416 234144 217508 234172
rect 136416 234132 136422 234144
rect 217502 234132 217508 234144
rect 217560 234132 217566 234184
rect 38838 234064 38844 234116
rect 38896 234104 38902 234116
rect 139394 234104 139400 234116
rect 38896 234076 139400 234104
rect 38896 234064 38902 234076
rect 139394 234064 139400 234076
rect 139452 234064 139458 234116
rect 170950 234064 170956 234116
rect 171008 234104 171014 234116
rect 217318 234104 217324 234116
rect 171008 234076 217324 234104
rect 171008 234064 171014 234076
rect 217318 234064 217324 234076
rect 217376 234064 217382 234116
rect 39022 233996 39028 234048
rect 39080 234036 39086 234048
rect 146294 234036 146300 234048
rect 39080 234008 146300 234036
rect 39080 233996 39086 234008
rect 146294 233996 146300 234008
rect 146352 233996 146358 234048
rect 150250 233996 150256 234048
rect 150308 234036 150314 234048
rect 247034 234036 247040 234048
rect 150308 234008 247040 234036
rect 150308 233996 150314 234008
rect 247034 233996 247040 234008
rect 247092 233996 247098 234048
rect 56502 233928 56508 233980
rect 56560 233968 56566 233980
rect 118234 233968 118240 233980
rect 56560 233940 118240 233968
rect 56560 233928 56566 233940
rect 118234 233928 118240 233940
rect 118292 233928 118298 233980
rect 129366 233928 129372 233980
rect 129424 233968 129430 233980
rect 235994 233968 236000 233980
rect 129424 233940 236000 233968
rect 129424 233928 129430 233940
rect 235994 233928 236000 233940
rect 236052 233928 236058 233980
rect 38286 233860 38292 233912
rect 38344 233900 38350 233912
rect 181070 233900 181076 233912
rect 38344 233872 181076 233900
rect 38344 233860 38350 233872
rect 181070 233860 181076 233872
rect 181128 233860 181134 233912
rect 77018 233044 77024 233096
rect 77076 233084 77082 233096
rect 142706 233084 142712 233096
rect 77076 233056 142712 233084
rect 77076 233044 77082 233056
rect 142706 233044 142712 233056
rect 142764 233044 142770 233096
rect 115382 232976 115388 233028
rect 115440 233016 115446 233028
rect 182818 233016 182824 233028
rect 115440 232988 182824 233016
rect 115440 232976 115446 232988
rect 182818 232976 182824 232988
rect 182876 232976 182882 233028
rect 185210 232976 185216 233028
rect 185268 233016 185274 233028
rect 202138 233016 202144 233028
rect 185268 232988 202144 233016
rect 185268 232976 185274 232988
rect 202138 232976 202144 232988
rect 202196 232976 202202 233028
rect 125870 232908 125876 232960
rect 125928 232948 125934 232960
rect 203518 232948 203524 232960
rect 125928 232920 203524 232948
rect 125928 232908 125934 232920
rect 203518 232908 203524 232920
rect 203576 232908 203582 232960
rect 213086 232908 213092 232960
rect 213144 232948 213150 232960
rect 284938 232948 284944 232960
rect 213144 232920 284944 232948
rect 213144 232908 213150 232920
rect 284938 232908 284944 232920
rect 284996 232908 285002 232960
rect 81250 232840 81256 232892
rect 81308 232880 81314 232892
rect 163590 232880 163596 232892
rect 81308 232852 163596 232880
rect 81308 232840 81314 232852
rect 163590 232840 163596 232852
rect 163648 232840 163654 232892
rect 202598 232840 202604 232892
rect 202656 232880 202662 232892
rect 282178 232880 282184 232892
rect 202656 232852 282184 232880
rect 202656 232840 202662 232852
rect 282178 232840 282184 232852
rect 282236 232840 282242 232892
rect 68830 232772 68836 232824
rect 68888 232812 68894 232824
rect 153194 232812 153200 232824
rect 68888 232784 153200 232812
rect 68888 232772 68894 232784
rect 153194 232772 153200 232784
rect 153252 232772 153258 232824
rect 162118 232772 162124 232824
rect 162176 232812 162182 232824
rect 258166 232812 258172 232824
rect 162176 232784 258172 232812
rect 162176 232772 162182 232784
rect 258166 232772 258172 232784
rect 258224 232772 258230 232824
rect 137278 232704 137284 232756
rect 137336 232744 137342 232756
rect 236822 232744 236828 232756
rect 137336 232716 236828 232744
rect 137336 232704 137342 232716
rect 236822 232704 236828 232716
rect 236880 232704 236886 232756
rect 242802 232704 242808 232756
rect 242860 232744 242866 232756
rect 261110 232744 261116 232756
rect 242860 232716 261116 232744
rect 242860 232704 242866 232716
rect 261110 232704 261116 232716
rect 261168 232704 261174 232756
rect 68738 232636 68744 232688
rect 68796 232676 68802 232688
rect 121730 232676 121736 232688
rect 68796 232648 121736 232676
rect 68796 232636 68802 232648
rect 121730 232636 121736 232648
rect 121788 232636 121794 232688
rect 140038 232636 140044 232688
rect 140096 232676 140102 232688
rect 247310 232676 247316 232688
rect 140096 232648 247316 232676
rect 140096 232636 140102 232648
rect 247310 232636 247316 232648
rect 247368 232636 247374 232688
rect 251082 232636 251088 232688
rect 251140 232676 251146 232688
rect 260834 232676 260840 232688
rect 251140 232648 260840 232676
rect 251140 232636 251146 232648
rect 260834 232636 260840 232648
rect 260892 232636 260898 232688
rect 111702 232568 111708 232620
rect 111760 232608 111766 232620
rect 219618 232608 219624 232620
rect 111760 232580 219624 232608
rect 111760 232568 111766 232580
rect 219618 232568 219624 232580
rect 219676 232568 219682 232620
rect 254946 232568 254952 232620
rect 255004 232608 255010 232620
rect 275278 232608 275284 232620
rect 255004 232580 275284 232608
rect 255004 232568 255010 232580
rect 275278 232568 275284 232580
rect 275336 232568 275342 232620
rect 114462 232500 114468 232552
rect 114520 232540 114526 232552
rect 226334 232540 226340 232552
rect 114520 232512 226340 232540
rect 114520 232500 114526 232512
rect 226334 232500 226340 232512
rect 226392 232500 226398 232552
rect 251450 232500 251456 232552
rect 251508 232540 251514 232552
rect 304258 232540 304264 232552
rect 251508 232512 304264 232540
rect 251508 232500 251514 232512
rect 304258 232500 304264 232512
rect 304316 232500 304322 232552
rect 217962 231752 217968 231804
rect 218020 231792 218026 231804
rect 262674 231792 262680 231804
rect 218020 231764 262680 231792
rect 218020 231752 218026 231764
rect 262674 231752 262680 231764
rect 262732 231752 262738 231804
rect 139302 231684 139308 231736
rect 139360 231724 139366 231736
rect 262950 231724 262956 231736
rect 139360 231696 262956 231724
rect 139360 231684 139366 231696
rect 262950 231684 262956 231696
rect 263008 231684 263014 231736
rect 133782 231616 133788 231668
rect 133840 231656 133846 231668
rect 262858 231656 262864 231668
rect 133840 231628 262864 231656
rect 133840 231616 133846 231628
rect 262858 231616 262864 231628
rect 262916 231616 262922 231668
rect 124122 231548 124128 231600
rect 124180 231588 124186 231600
rect 262766 231588 262772 231600
rect 124180 231560 262772 231588
rect 124180 231548 124186 231560
rect 262766 231548 262772 231560
rect 262824 231548 262830 231600
rect 109494 231480 109500 231532
rect 109552 231520 109558 231532
rect 115934 231520 115940 231532
rect 109552 231492 115940 231520
rect 109552 231480 109558 231492
rect 115934 231480 115940 231492
rect 115992 231480 115998 231532
rect 121362 231480 121368 231532
rect 121420 231520 121426 231532
rect 261294 231520 261300 231532
rect 121420 231492 261300 231520
rect 121420 231480 121426 231492
rect 261294 231480 261300 231492
rect 261352 231480 261358 231532
rect 108206 231412 108212 231464
rect 108264 231452 108270 231464
rect 252554 231452 252560 231464
rect 108264 231424 252560 231452
rect 108264 231412 108270 231424
rect 252554 231412 252560 231424
rect 252612 231412 252618 231464
rect 256602 231412 256608 231464
rect 256660 231452 256666 231464
rect 261202 231452 261208 231464
rect 256660 231424 261208 231452
rect 256660 231412 256666 231424
rect 261202 231412 261208 231424
rect 261260 231412 261266 231464
rect 108298 231344 108304 231396
rect 108356 231384 108362 231396
rect 258074 231384 258080 231396
rect 108356 231356 258080 231384
rect 108356 231344 108362 231356
rect 258074 231344 258080 231356
rect 258132 231344 258138 231396
rect 91002 231276 91008 231328
rect 91060 231316 91066 231328
rect 262398 231316 262404 231328
rect 91060 231288 262404 231316
rect 91060 231276 91066 231288
rect 262398 231276 262404 231288
rect 262456 231276 262462 231328
rect 108482 231208 108488 231260
rect 108540 231248 108546 231260
rect 322934 231248 322940 231260
rect 108540 231220 322940 231248
rect 108540 231208 108546 231220
rect 322934 231208 322940 231220
rect 322992 231208 322998 231260
rect 60550 231140 60556 231192
rect 60608 231180 60614 231192
rect 261018 231180 261024 231192
rect 60608 231152 261024 231180
rect 60608 231140 60614 231152
rect 261018 231140 261024 231152
rect 261076 231140 261082 231192
rect 110322 231072 110328 231124
rect 110380 231112 110386 231124
rect 325694 231112 325700 231124
rect 110380 231084 325700 231112
rect 110380 231072 110386 231084
rect 325694 231072 325700 231084
rect 325752 231072 325758 231124
rect 237282 231004 237288 231056
rect 237340 231044 237346 231056
rect 260466 231044 260472 231056
rect 237340 231016 260472 231044
rect 237340 231004 237346 231016
rect 260466 231004 260472 231016
rect 260524 231004 260530 231056
rect 240042 230936 240048 230988
rect 240100 230976 240106 230988
rect 260558 230976 260564 230988
rect 240100 230948 260564 230976
rect 240100 230936 240106 230948
rect 260558 230936 260564 230948
rect 260616 230936 260622 230988
rect 146202 230392 146208 230444
rect 146260 230432 146266 230444
rect 259362 230432 259368 230444
rect 146260 230404 259368 230432
rect 146260 230392 146266 230404
rect 259362 230392 259368 230404
rect 259420 230392 259426 230444
rect 217870 230052 217876 230104
rect 217928 230092 217934 230104
rect 263042 230092 263048 230104
rect 217928 230064 263048 230092
rect 217928 230052 217934 230064
rect 263042 230052 263048 230064
rect 263100 230052 263106 230104
rect 248322 229984 248328 230036
rect 248380 230024 248386 230036
rect 260006 230024 260012 230036
rect 248380 229996 260012 230024
rect 248380 229984 248386 229996
rect 260006 229984 260012 229996
rect 260064 229984 260070 230036
rect 99190 229916 99196 229968
rect 99248 229956 99254 229968
rect 259914 229956 259920 229968
rect 99248 229928 259920 229956
rect 99248 229916 99254 229928
rect 259914 229916 259920 229928
rect 259972 229916 259978 229968
rect 108390 229848 108396 229900
rect 108448 229888 108454 229900
rect 262582 229888 262588 229900
rect 108448 229860 262588 229888
rect 108448 229848 108454 229860
rect 262582 229848 262588 229860
rect 262640 229848 262646 229900
rect 99098 229780 99104 229832
rect 99156 229820 99162 229832
rect 259822 229820 259828 229832
rect 99156 229792 259828 229820
rect 99156 229780 99162 229792
rect 259822 229780 259828 229792
rect 259880 229780 259886 229832
rect 96430 229712 96436 229764
rect 96488 229752 96494 229764
rect 262490 229752 262496 229764
rect 96488 229724 262496 229752
rect 96488 229712 96494 229724
rect 262490 229712 262496 229724
rect 262548 229712 262554 229764
rect 263502 224884 263508 224936
rect 263560 224924 263566 224936
rect 276658 224924 276664 224936
rect 263560 224896 276664 224924
rect 263560 224884 263566 224896
rect 276658 224884 276664 224896
rect 276716 224884 276722 224936
rect 261110 224272 261116 224324
rect 261168 224272 261174 224324
rect 259822 224204 259828 224256
rect 259880 224244 259886 224256
rect 260466 224244 260472 224256
rect 259880 224216 260472 224244
rect 259880 224204 259886 224216
rect 260466 224204 260472 224216
rect 260524 224204 260530 224256
rect 261128 224120 261156 224272
rect 262306 224204 262312 224256
rect 262364 224244 262370 224256
rect 262674 224244 262680 224256
rect 262364 224216 262680 224244
rect 262364 224204 262370 224216
rect 262674 224204 262680 224216
rect 262732 224204 262738 224256
rect 261110 224068 261116 224120
rect 261168 224068 261174 224120
rect 262766 223864 262772 223916
rect 262824 223864 262830 223916
rect 262784 223712 262812 223864
rect 262766 223660 262772 223712
rect 262824 223660 262830 223712
rect 97902 223524 97908 223576
rect 97960 223564 97966 223576
rect 107654 223564 107660 223576
rect 97960 223536 107660 223564
rect 97960 223524 97966 223536
rect 107654 223524 107660 223536
rect 107712 223524 107718 223576
rect 262950 223524 262956 223576
rect 263008 223564 263014 223576
rect 305638 223564 305644 223576
rect 263008 223536 305644 223564
rect 263008 223524 263014 223536
rect 305638 223524 305644 223536
rect 305696 223524 305702 223576
rect 260006 222164 260012 222216
rect 260064 222204 260070 222216
rect 260558 222204 260564 222216
rect 260064 222176 260564 222204
rect 260064 222164 260070 222176
rect 260558 222164 260564 222176
rect 260616 222164 260622 222216
rect 93670 217948 93676 218000
rect 93728 217988 93734 218000
rect 107654 217988 107660 218000
rect 93728 217960 107660 217988
rect 93728 217948 93734 217960
rect 107654 217948 107660 217960
rect 107712 217948 107718 218000
rect 263502 217948 263508 218000
rect 263560 217988 263566 218000
rect 300118 217988 300124 218000
rect 263560 217960 300124 217988
rect 263560 217948 263566 217960
rect 300118 217948 300124 217960
rect 300176 217948 300182 218000
rect 263502 216588 263508 216640
rect 263560 216628 263566 216640
rect 298738 216628 298744 216640
rect 263560 216600 298744 216628
rect 263560 216588 263566 216600
rect 298738 216588 298744 216600
rect 298796 216588 298802 216640
rect 263502 213868 263508 213920
rect 263560 213908 263566 213920
rect 294598 213908 294604 213920
rect 263560 213880 294604 213908
rect 263560 213868 263566 213880
rect 294598 213868 294604 213880
rect 294656 213868 294662 213920
rect 263502 211080 263508 211132
rect 263560 211120 263566 211132
rect 291838 211120 291844 211132
rect 263560 211092 291844 211120
rect 263560 211080 263566 211092
rect 291838 211080 291844 211092
rect 291896 211080 291902 211132
rect 263502 204212 263508 204264
rect 263560 204252 263566 204264
rect 277486 204252 277492 204264
rect 263560 204224 277492 204252
rect 263560 204212 263566 204224
rect 277486 204212 277492 204224
rect 277544 204212 277550 204264
rect 262214 189932 262220 189984
rect 262272 189972 262278 189984
rect 264330 189972 264336 189984
rect 262272 189944 264336 189972
rect 262272 189932 262278 189944
rect 264330 189932 264336 189944
rect 264388 189932 264394 189984
rect 75822 188980 75828 189032
rect 75880 189020 75886 189032
rect 107654 189020 107660 189032
rect 75880 188992 107660 189020
rect 75880 188980 75886 188992
rect 107654 188980 107660 188992
rect 107712 188980 107718 189032
rect 88150 186260 88156 186312
rect 88208 186300 88214 186312
rect 107654 186300 107660 186312
rect 88208 186272 107660 186300
rect 88208 186260 88214 186272
rect 107654 186260 107660 186272
rect 107712 186260 107718 186312
rect 38746 180752 38752 180804
rect 38804 180792 38810 180804
rect 107654 180792 107660 180804
rect 38804 180764 107660 180792
rect 38804 180752 38810 180764
rect 107654 180752 107660 180764
rect 107712 180752 107718 180804
rect 78490 177964 78496 178016
rect 78548 178004 78554 178016
rect 107654 178004 107660 178016
rect 78548 177976 107660 178004
rect 78548 177964 78554 177976
rect 107654 177964 107660 177976
rect 107712 177964 107718 178016
rect 62022 172456 62028 172508
rect 62080 172496 62086 172508
rect 107654 172496 107660 172508
rect 62080 172468 107660 172496
rect 62080 172456 62086 172468
rect 107654 172456 107660 172468
rect 107712 172456 107718 172508
rect 74442 169668 74448 169720
rect 74500 169708 74506 169720
rect 107654 169708 107660 169720
rect 74500 169680 107660 169708
rect 74500 169668 74506 169680
rect 107654 169668 107660 169680
rect 107712 169668 107718 169720
rect 63402 164160 63408 164212
rect 63460 164200 63466 164212
rect 107654 164200 107660 164212
rect 63460 164172 107660 164200
rect 63460 164160 63466 164172
rect 107654 164160 107660 164172
rect 107712 164160 107718 164212
rect 38470 161372 38476 161424
rect 38528 161412 38534 161424
rect 107654 161412 107660 161424
rect 38528 161384 107660 161412
rect 38528 161372 38534 161384
rect 107654 161372 107660 161384
rect 107712 161372 107718 161424
rect 96522 160420 96528 160472
rect 96580 160460 96586 160472
rect 110598 160460 110604 160472
rect 96580 160432 110604 160460
rect 96580 160420 96586 160432
rect 110598 160420 110604 160432
rect 110656 160420 110662 160472
rect 260374 160080 260380 160132
rect 260432 160120 260438 160132
rect 263686 160120 263692 160132
rect 260432 160092 263692 160120
rect 260432 160080 260438 160092
rect 263686 160080 263692 160092
rect 263744 160080 263750 160132
rect 242802 159400 242808 159452
rect 242860 159440 242866 159452
rect 273346 159440 273352 159452
rect 242860 159412 273352 159440
rect 242860 159400 242866 159412
rect 273346 159400 273352 159412
rect 273404 159400 273410 159452
rect 110414 159332 110420 159384
rect 110472 159372 110478 159384
rect 111150 159372 111156 159384
rect 110472 159344 111156 159372
rect 110472 159332 110478 159344
rect 111150 159332 111156 159344
rect 111208 159332 111214 159384
rect 244274 159332 244280 159384
rect 244332 159372 244338 159384
rect 282914 159372 282920 159384
rect 244332 159344 282920 159372
rect 244332 159332 244338 159344
rect 282914 159332 282920 159344
rect 282972 159332 282978 159384
rect 85482 159264 85488 159316
rect 85540 159304 85546 159316
rect 240686 159304 240692 159316
rect 85540 159276 240692 159304
rect 85540 159264 85546 159276
rect 240686 159264 240692 159276
rect 240744 159264 240750 159316
rect 78582 159196 78588 159248
rect 78640 159236 78646 159248
rect 233510 159236 233516 159248
rect 78640 159208 233516 159236
rect 78640 159196 78646 159208
rect 233510 159196 233516 159208
rect 233568 159196 233574 159248
rect 256602 159196 256608 159248
rect 256660 159236 256666 159248
rect 274634 159236 274640 159248
rect 256660 159208 274640 159236
rect 256660 159196 256666 159208
rect 274634 159196 274640 159208
rect 274692 159196 274698 159248
rect 86770 159128 86776 159180
rect 86828 159168 86834 159180
rect 243722 159168 243728 159180
rect 86828 159140 243728 159168
rect 86828 159128 86834 159140
rect 243722 159128 243728 159140
rect 243780 159128 243786 159180
rect 246390 159128 246396 159180
rect 246448 159168 246454 159180
rect 266446 159168 266452 159180
rect 246448 159140 266452 159168
rect 246448 159128 246454 159140
rect 266446 159128 266452 159140
rect 266504 159128 266510 159180
rect 92290 159060 92296 159112
rect 92348 159100 92354 159112
rect 249886 159100 249892 159112
rect 92348 159072 249892 159100
rect 92348 159060 92354 159072
rect 249886 159060 249892 159072
rect 249944 159060 249950 159112
rect 253566 159060 253572 159112
rect 253624 159100 253630 159112
rect 273254 159100 273260 159112
rect 253624 159072 273260 159100
rect 253624 159060 253630 159072
rect 273254 159060 273260 159072
rect 273312 159060 273318 159112
rect 95142 158992 95148 159044
rect 95200 159032 95206 159044
rect 253934 159032 253940 159044
rect 95200 159004 253940 159032
rect 95200 158992 95206 159004
rect 253934 158992 253940 159004
rect 253992 158992 253998 159044
rect 259362 158992 259368 159044
rect 259420 159032 259426 159044
rect 278774 159032 278780 159044
rect 259420 159004 278780 159032
rect 259420 158992 259426 159004
rect 278774 158992 278780 159004
rect 278832 158992 278838 159044
rect 88242 158924 88248 158976
rect 88300 158964 88306 158976
rect 247126 158964 247132 158976
rect 88300 158936 247132 158964
rect 88300 158924 88306 158936
rect 247126 158924 247132 158936
rect 247184 158924 247190 158976
rect 249518 158924 249524 158976
rect 249576 158964 249582 158976
rect 270586 158964 270592 158976
rect 249576 158936 270592 158964
rect 249576 158924 249582 158936
rect 270586 158924 270592 158936
rect 270644 158924 270650 158976
rect 38654 158856 38660 158908
rect 38712 158896 38718 158908
rect 217226 158896 217232 158908
rect 38712 158868 217232 158896
rect 38712 158856 38718 158868
rect 217226 158856 217232 158868
rect 217284 158856 217290 158908
rect 243354 158856 243360 158908
rect 243412 158896 243418 158908
rect 266354 158896 266360 158908
rect 243412 158868 266360 158896
rect 243412 158856 243418 158868
rect 266354 158856 266360 158868
rect 266412 158856 266418 158908
rect 38562 158788 38568 158840
rect 38620 158828 38626 158840
rect 224310 158828 224316 158840
rect 38620 158800 224316 158828
rect 38620 158788 38626 158800
rect 224310 158788 224316 158800
rect 224368 158788 224374 158840
rect 240042 158788 240048 158840
rect 240100 158828 240106 158840
rect 263594 158828 263600 158840
rect 240100 158800 263600 158828
rect 240100 158788 240106 158800
rect 263594 158788 263600 158800
rect 263652 158788 263658 158840
rect 39942 158720 39948 158772
rect 40000 158760 40006 158772
rect 110414 158760 110420 158772
rect 40000 158732 110420 158760
rect 40000 158720 40006 158732
rect 110414 158720 110420 158732
rect 110472 158720 110478 158772
rect 113174 158720 113180 158772
rect 113232 158760 113238 158772
rect 383654 158760 383660 158772
rect 113232 158732 383660 158760
rect 113232 158720 113238 158732
rect 383654 158720 383660 158732
rect 383712 158720 383718 158772
rect 60642 158652 60648 158704
rect 60700 158692 60706 158704
rect 219434 158692 219440 158704
rect 60700 158664 219440 158692
rect 60700 158652 60706 158664
rect 219434 158652 219440 158664
rect 219492 158652 219498 158704
rect 235902 158652 235908 158704
rect 235960 158692 235966 158704
rect 244274 158692 244280 158704
rect 235960 158664 244280 158692
rect 235960 158652 235966 158664
rect 244274 158652 244280 158664
rect 244332 158652 244338 158704
rect 248230 158652 248236 158704
rect 248288 158692 248294 158704
rect 295978 158692 295984 158704
rect 248288 158664 295984 158692
rect 248288 158652 248294 158664
rect 295978 158652 295984 158664
rect 296036 158652 296042 158704
rect 92382 158584 92388 158636
rect 92440 158624 92446 158636
rect 251266 158624 251272 158636
rect 92440 158596 251272 158624
rect 92440 158584 92446 158596
rect 251266 158584 251272 158596
rect 251324 158584 251330 158636
rect 255590 158584 255596 158636
rect 255648 158624 255654 158636
rect 302878 158624 302884 158636
rect 255648 158596 302884 158624
rect 255648 158584 255654 158596
rect 302878 158584 302884 158596
rect 302936 158584 302942 158636
rect 69658 158516 69664 158568
rect 69716 158556 69722 158568
rect 225322 158556 225328 158568
rect 69716 158528 225328 158556
rect 69716 158516 69722 158528
rect 225322 158516 225328 158528
rect 225380 158516 225386 158568
rect 239306 158516 239312 158568
rect 239364 158556 239370 158568
rect 286318 158556 286324 158568
rect 239364 158528 286324 158556
rect 239364 158516 239370 158528
rect 286318 158516 286324 158528
rect 286376 158516 286382 158568
rect 59262 158448 59268 158500
rect 59320 158488 59326 158500
rect 214190 158488 214196 158500
rect 59320 158460 214196 158488
rect 59320 158448 59326 158460
rect 214190 158448 214196 158460
rect 214248 158448 214254 158500
rect 242342 158448 242348 158500
rect 242400 158488 242406 158500
rect 287698 158488 287704 158500
rect 242400 158460 287704 158488
rect 242400 158448 242406 158460
rect 287698 158448 287704 158460
rect 287756 158448 287762 158500
rect 67542 158380 67548 158432
rect 67600 158420 67606 158432
rect 221274 158420 221280 158432
rect 67600 158392 221280 158420
rect 67600 158380 67606 158392
rect 221274 158380 221280 158392
rect 221332 158380 221338 158432
rect 231118 158380 231124 158432
rect 231176 158420 231182 158432
rect 242802 158420 242808 158432
rect 231176 158392 242808 158420
rect 231176 158380 231182 158392
rect 242802 158380 242808 158392
rect 242860 158380 242866 158432
rect 245378 158380 245384 158432
rect 245436 158420 245442 158432
rect 289078 158420 289084 158432
rect 245436 158392 289084 158420
rect 245436 158380 245442 158392
rect 289078 158380 289084 158392
rect 289136 158380 289142 158432
rect 110598 158312 110604 158364
rect 110656 158352 110662 158364
rect 256970 158352 256976 158364
rect 110656 158324 256976 158352
rect 110656 158312 110662 158324
rect 256970 158312 256976 158324
rect 257028 158312 257034 158364
rect 230106 158244 230112 158296
rect 230164 158284 230170 158296
rect 270494 158284 270500 158296
rect 230164 158256 270500 158284
rect 230164 158244 230170 158256
rect 270494 158244 270500 158256
rect 270552 158244 270558 158296
rect 227070 158176 227076 158228
rect 227128 158216 227134 158228
rect 260374 158216 260380 158228
rect 227128 158188 260380 158216
rect 227128 158176 227134 158188
rect 260374 158176 260380 158188
rect 260432 158176 260438 158228
rect 102042 158108 102048 158160
rect 102100 158148 102106 158160
rect 234614 158148 234620 158160
rect 102100 158120 234620 158148
rect 102100 158108 102106 158120
rect 234614 158108 234620 158120
rect 234672 158108 234678 158160
rect 104802 158040 104808 158092
rect 104860 158080 104866 158092
rect 236546 158080 236552 158092
rect 104860 158052 236552 158080
rect 104860 158040 104866 158052
rect 236546 158040 236552 158052
rect 236604 158040 236610 158092
rect 106182 157972 106188 158024
rect 106240 158012 106246 158024
rect 237650 158012 237656 158024
rect 106240 157984 237656 158012
rect 106240 157972 106246 157984
rect 237650 157972 237656 157984
rect 237708 157972 237714 158024
rect 228082 157904 228088 157956
rect 228140 157944 228146 157956
rect 264238 157944 264244 157956
rect 228140 157916 264244 157944
rect 228140 157904 228146 157916
rect 264238 157904 264244 157916
rect 264296 157904 264302 157956
rect 99282 157836 99288 157888
rect 99340 157876 99346 157888
rect 232498 157876 232504 157888
rect 99340 157848 232504 157876
rect 99340 157836 99346 157848
rect 232498 157836 232504 157848
rect 232556 157836 232562 157888
rect 93762 157768 93768 157820
rect 93820 157808 93826 157820
rect 231854 157808 231860 157820
rect 93820 157780 231860 157808
rect 93820 157768 93826 157780
rect 231854 157768 231860 157780
rect 231912 157768 231918 157820
rect 114554 155932 114560 155984
rect 114612 155972 114618 155984
rect 115198 155972 115204 155984
rect 114612 155944 115204 155972
rect 114612 155932 114618 155944
rect 115198 155932 115204 155944
rect 115256 155932 115262 155984
rect 117314 155932 117320 155984
rect 117372 155972 117378 155984
rect 118234 155972 118240 155984
rect 117372 155944 118240 155972
rect 117372 155932 117378 155944
rect 118234 155932 118240 155944
rect 118292 155932 118298 155984
rect 121454 155932 121460 155984
rect 121512 155972 121518 155984
rect 122374 155972 122380 155984
rect 121512 155944 122380 155972
rect 121512 155932 121518 155944
rect 122374 155932 122380 155944
rect 122432 155932 122438 155984
rect 129734 155932 129740 155984
rect 129792 155972 129798 155984
rect 130470 155972 130476 155984
rect 129792 155944 130476 155972
rect 129792 155932 129798 155944
rect 130470 155932 130476 155944
rect 130528 155932 130534 155984
rect 133874 155932 133880 155984
rect 133932 155972 133938 155984
rect 134610 155972 134616 155984
rect 133932 155944 134616 155972
rect 133932 155932 133938 155944
rect 134610 155932 134616 155944
rect 134668 155932 134674 155984
rect 144914 155932 144920 155984
rect 144972 155972 144978 155984
rect 145834 155972 145840 155984
rect 144972 155944 145840 155972
rect 144972 155932 144978 155944
rect 145834 155932 145840 155944
rect 145892 155932 145898 155984
rect 149054 155932 149060 155984
rect 149112 155972 149118 155984
rect 149882 155972 149888 155984
rect 149112 155944 149888 155972
rect 149112 155932 149118 155944
rect 149882 155932 149888 155944
rect 149940 155932 149946 155984
rect 157334 155932 157340 155984
rect 157392 155972 157398 155984
rect 158070 155972 158076 155984
rect 157392 155944 158076 155972
rect 157392 155932 157398 155944
rect 158070 155932 158076 155944
rect 158128 155932 158134 155984
rect 161474 155932 161480 155984
rect 161532 155972 161538 155984
rect 162118 155972 162124 155984
rect 161532 155944 162124 155972
rect 161532 155932 161538 155944
rect 162118 155932 162124 155944
rect 162176 155932 162182 155984
rect 164234 155932 164240 155984
rect 164292 155972 164298 155984
rect 165154 155972 165160 155984
rect 164292 155944 165160 155972
rect 164292 155932 164298 155944
rect 165154 155932 165160 155944
rect 165212 155932 165218 155984
rect 172514 155932 172520 155984
rect 172572 155972 172578 155984
rect 173342 155972 173348 155984
rect 172572 155944 173348 155972
rect 172572 155932 172578 155944
rect 173342 155932 173348 155944
rect 173400 155932 173406 155984
rect 176654 155932 176660 155984
rect 176712 155972 176718 155984
rect 177390 155972 177396 155984
rect 176712 155944 177396 155972
rect 176712 155932 176718 155944
rect 177390 155932 177396 155944
rect 177448 155932 177454 155984
rect 184934 155932 184940 155984
rect 184992 155972 184998 155984
rect 185578 155972 185584 155984
rect 184992 155944 185584 155972
rect 184992 155932 184998 155944
rect 185578 155932 185584 155944
rect 185636 155932 185642 155984
rect 187694 155932 187700 155984
rect 187752 155972 187758 155984
rect 188614 155972 188620 155984
rect 187752 155944 188620 155972
rect 187752 155932 187758 155944
rect 188614 155932 188620 155944
rect 188672 155932 188678 155984
rect 200114 155932 200120 155984
rect 200172 155972 200178 155984
rect 200850 155972 200856 155984
rect 200172 155944 200856 155972
rect 200172 155932 200178 155944
rect 200850 155932 200856 155944
rect 200908 155932 200914 155984
rect 204254 155932 204260 155984
rect 204312 155972 204318 155984
rect 204990 155972 204996 155984
rect 204312 155944 204996 155972
rect 204312 155932 204318 155944
rect 204990 155932 204996 155944
rect 205048 155932 205054 155984
rect 191834 153688 191840 153740
rect 191892 153728 191898 153740
rect 192754 153728 192760 153740
rect 191892 153700 192760 153728
rect 191892 153688 191898 153700
rect 192754 153688 192760 153700
rect 192812 153688 192818 153740
rect 111794 120028 111800 120080
rect 111852 120068 111858 120080
rect 256694 120068 256700 120080
rect 111852 120040 256700 120068
rect 111852 120028 111858 120040
rect 256694 120028 256700 120040
rect 256752 120028 256758 120080
rect 342254 120028 342260 120080
rect 342312 120068 342318 120080
rect 382274 120068 382280 120080
rect 342312 120040 382280 120068
rect 342312 120028 342318 120040
rect 382274 120028 382280 120040
rect 382332 120028 382338 120080
rect 110506 118600 110512 118652
rect 110564 118640 110570 118652
rect 256694 118640 256700 118652
rect 110564 118612 256700 118640
rect 110564 118600 110570 118612
rect 256694 118600 256700 118612
rect 256752 118600 256758 118652
rect 342346 118600 342352 118652
rect 342404 118640 342410 118652
rect 386414 118640 386420 118652
rect 342404 118612 386420 118640
rect 342404 118600 342410 118612
rect 386414 118600 386420 118612
rect 386472 118600 386478 118652
rect 114646 118532 114652 118584
rect 114704 118572 114710 118584
rect 256786 118572 256792 118584
rect 114704 118544 256792 118572
rect 114704 118532 114710 118544
rect 256786 118532 256792 118544
rect 256844 118532 256850 118584
rect 342254 118532 342260 118584
rect 342312 118572 342318 118584
rect 379514 118572 379520 118584
rect 342312 118544 379520 118572
rect 342312 118532 342318 118544
rect 379514 118532 379520 118544
rect 379572 118532 379578 118584
rect 114554 117240 114560 117292
rect 114612 117280 114618 117292
rect 256694 117280 256700 117292
rect 114612 117252 256700 117280
rect 114612 117240 114618 117252
rect 256694 117240 256700 117252
rect 256752 117240 256758 117292
rect 342346 117240 342352 117292
rect 342404 117280 342410 117292
rect 518158 117280 518164 117292
rect 342404 117252 518164 117280
rect 342404 117240 342410 117252
rect 518158 117240 518164 117252
rect 518216 117240 518222 117292
rect 211246 117172 211252 117224
rect 211304 117212 211310 117224
rect 256786 117212 256792 117224
rect 211304 117184 256792 117212
rect 211304 117172 211310 117184
rect 256786 117172 256792 117184
rect 256844 117172 256850 117224
rect 342254 117172 342260 117224
rect 342312 117212 342318 117224
rect 387794 117212 387800 117224
rect 342312 117184 387800 117212
rect 342312 117172 342318 117184
rect 387794 117172 387800 117184
rect 387852 117172 387858 117224
rect 205634 115880 205640 115932
rect 205692 115920 205698 115932
rect 256786 115920 256792 115932
rect 205692 115892 256792 115920
rect 205692 115880 205698 115892
rect 256786 115880 256792 115892
rect 256844 115880 256850 115932
rect 342254 115880 342260 115932
rect 342312 115920 342318 115932
rect 512638 115920 512644 115932
rect 342312 115892 512644 115920
rect 342312 115880 342318 115892
rect 512638 115880 512644 115892
rect 512696 115880 512702 115932
rect 208486 115812 208492 115864
rect 208544 115852 208550 115864
rect 256694 115852 256700 115864
rect 208544 115824 256700 115852
rect 208544 115812 208550 115824
rect 256694 115812 256700 115824
rect 256752 115812 256758 115864
rect 342346 115812 342352 115864
rect 342404 115852 342410 115864
rect 508498 115852 508504 115864
rect 342404 115824 508504 115852
rect 342404 115812 342410 115824
rect 508498 115812 508504 115824
rect 508556 115812 508562 115864
rect 202874 114452 202880 114504
rect 202932 114492 202938 114504
rect 256694 114492 256700 114504
rect 202932 114464 256700 114492
rect 202932 114452 202938 114464
rect 256694 114452 256700 114464
rect 256752 114452 256758 114504
rect 342254 114452 342260 114504
rect 342312 114492 342318 114504
rect 504358 114492 504364 114504
rect 342312 114464 504364 114492
rect 342312 114452 342318 114464
rect 504358 114452 504364 114464
rect 504416 114452 504422 114504
rect 196066 113092 196072 113144
rect 196124 113132 196130 113144
rect 256786 113132 256792 113144
rect 196124 113104 256792 113132
rect 196124 113092 196130 113104
rect 256786 113092 256792 113104
rect 256844 113092 256850 113144
rect 342254 113092 342260 113144
rect 342312 113132 342318 113144
rect 501598 113132 501604 113144
rect 342312 113104 501604 113132
rect 342312 113092 342318 113104
rect 501598 113092 501604 113104
rect 501656 113092 501662 113144
rect 200206 113024 200212 113076
rect 200264 113064 200270 113076
rect 256694 113064 256700 113076
rect 200264 113036 256700 113064
rect 200264 113024 200270 113036
rect 256694 113024 256700 113036
rect 256752 113024 256758 113076
rect 342346 113024 342352 113076
rect 342404 113064 342410 113076
rect 500218 113064 500224 113076
rect 342404 113036 500224 113064
rect 342404 113024 342410 113036
rect 500218 113024 500224 113036
rect 500276 113024 500282 113076
rect 190454 111732 190460 111784
rect 190512 111772 190518 111784
rect 256786 111772 256792 111784
rect 190512 111744 256792 111772
rect 190512 111732 190518 111744
rect 256786 111732 256792 111744
rect 256844 111732 256850 111784
rect 342254 111732 342260 111784
rect 342312 111772 342318 111784
rect 497458 111772 497464 111784
rect 342312 111744 497464 111772
rect 342312 111732 342318 111744
rect 497458 111732 497464 111744
rect 497516 111732 497522 111784
rect 193214 111664 193220 111716
rect 193272 111704 193278 111716
rect 256694 111704 256700 111716
rect 193272 111676 256700 111704
rect 193272 111664 193278 111676
rect 256694 111664 256700 111676
rect 256752 111664 256758 111716
rect 342346 111664 342352 111716
rect 342404 111704 342410 111716
rect 494698 111704 494704 111716
rect 342404 111676 494704 111704
rect 342404 111664 342410 111676
rect 494698 111664 494704 111676
rect 494756 111664 494762 111716
rect 187786 110372 187792 110424
rect 187844 110412 187850 110424
rect 256694 110412 256700 110424
rect 187844 110384 256700 110412
rect 187844 110372 187850 110384
rect 256694 110372 256700 110384
rect 256752 110372 256758 110424
rect 342254 110372 342260 110424
rect 342312 110412 342318 110424
rect 490558 110412 490564 110424
rect 342312 110384 490564 110412
rect 342312 110372 342318 110384
rect 490558 110372 490564 110384
rect 490616 110372 490622 110424
rect 180886 108944 180892 108996
rect 180944 108984 180950 108996
rect 256786 108984 256792 108996
rect 180944 108956 256792 108984
rect 180944 108944 180950 108956
rect 256786 108944 256792 108956
rect 256844 108944 256850 108996
rect 342254 108944 342260 108996
rect 342312 108984 342318 108996
rect 486418 108984 486424 108996
rect 342312 108956 486424 108984
rect 342312 108944 342318 108956
rect 486418 108944 486424 108956
rect 486476 108944 486482 108996
rect 185026 108876 185032 108928
rect 185084 108916 185090 108928
rect 256694 108916 256700 108928
rect 185084 108888 256700 108916
rect 185084 108876 185090 108888
rect 256694 108876 256700 108888
rect 256752 108876 256758 108928
rect 342346 108876 342352 108928
rect 342404 108916 342410 108928
rect 483014 108916 483020 108928
rect 342404 108888 483020 108916
rect 342404 108876 342410 108888
rect 483014 108876 483020 108888
rect 483072 108876 483078 108928
rect 175274 107584 175280 107636
rect 175332 107624 175338 107636
rect 256786 107624 256792 107636
rect 175332 107596 256792 107624
rect 175332 107584 175338 107596
rect 256786 107584 256792 107596
rect 256844 107584 256850 107636
rect 342254 107584 342260 107636
rect 342312 107624 342318 107636
rect 478874 107624 478880 107636
rect 342312 107596 478880 107624
rect 342312 107584 342318 107596
rect 478874 107584 478880 107596
rect 478932 107584 478938 107636
rect 178034 107516 178040 107568
rect 178092 107556 178098 107568
rect 256694 107556 256700 107568
rect 178092 107528 256700 107556
rect 178092 107516 178098 107528
rect 256694 107516 256700 107528
rect 256752 107516 256758 107568
rect 342346 107516 342352 107568
rect 342404 107556 342410 107568
rect 393958 107556 393964 107568
rect 342404 107528 393964 107556
rect 342404 107516 342410 107528
rect 393958 107516 393964 107528
rect 394016 107516 394022 107568
rect 168466 106224 168472 106276
rect 168524 106264 168530 106276
rect 256786 106264 256792 106276
rect 168524 106236 256792 106264
rect 168524 106224 168530 106236
rect 256786 106224 256792 106236
rect 256844 106224 256850 106276
rect 342346 106224 342352 106276
rect 342404 106264 342410 106276
rect 465074 106264 465080 106276
rect 342404 106236 465080 106264
rect 342404 106224 342410 106236
rect 465074 106224 465080 106236
rect 465132 106224 465138 106276
rect 172606 106156 172612 106208
rect 172664 106196 172670 106208
rect 256694 106196 256700 106208
rect 172664 106168 256700 106196
rect 172664 106156 172670 106168
rect 256694 106156 256700 106168
rect 256752 106156 256758 106208
rect 342254 106156 342260 106208
rect 342312 106196 342318 106208
rect 392578 106196 392584 106208
rect 342312 106168 392584 106196
rect 342312 106156 342318 106168
rect 392578 106156 392584 106168
rect 392636 106156 392642 106208
rect 165614 104796 165620 104848
rect 165672 104836 165678 104848
rect 256694 104836 256700 104848
rect 165672 104808 256700 104836
rect 165672 104796 165678 104808
rect 256694 104796 256700 104808
rect 256752 104796 256758 104848
rect 342254 104796 342260 104848
rect 342312 104836 342318 104848
rect 460934 104836 460940 104848
rect 342312 104808 460940 104836
rect 342312 104796 342318 104808
rect 460934 104796 460940 104808
rect 460992 104796 460998 104848
rect 160094 103436 160100 103488
rect 160152 103476 160158 103488
rect 256786 103476 256792 103488
rect 160152 103448 256792 103476
rect 160152 103436 160158 103448
rect 256786 103436 256792 103448
rect 256844 103436 256850 103488
rect 342254 103436 342260 103488
rect 342312 103476 342318 103488
rect 456794 103476 456800 103488
rect 342312 103448 456800 103476
rect 342312 103436 342318 103448
rect 456794 103436 456800 103448
rect 456852 103436 456858 103488
rect 162854 103368 162860 103420
rect 162912 103408 162918 103420
rect 256694 103408 256700 103420
rect 162912 103380 256700 103408
rect 162912 103368 162918 103380
rect 256694 103368 256700 103380
rect 256752 103368 256758 103420
rect 342346 103368 342352 103420
rect 342404 103408 342410 103420
rect 452654 103408 452660 103420
rect 342404 103380 452660 103408
rect 342404 103368 342410 103380
rect 452654 103368 452660 103380
rect 452712 103368 452718 103420
rect 153286 102076 153292 102128
rect 153344 102116 153350 102128
rect 256786 102116 256792 102128
rect 153344 102088 256792 102116
rect 153344 102076 153350 102088
rect 256786 102076 256792 102088
rect 256844 102076 256850 102128
rect 342254 102076 342260 102128
rect 342312 102116 342318 102128
rect 447134 102116 447140 102128
rect 342312 102088 447140 102116
rect 342312 102076 342318 102088
rect 447134 102076 447140 102088
rect 447192 102076 447198 102128
rect 157426 102008 157432 102060
rect 157484 102048 157490 102060
rect 256694 102048 256700 102060
rect 157484 102020 256700 102048
rect 157484 102008 157490 102020
rect 256694 102008 256700 102020
rect 256752 102008 256758 102060
rect 342346 102008 342352 102060
rect 342404 102048 342410 102060
rect 442994 102048 443000 102060
rect 342404 102020 443000 102048
rect 342404 102008 342410 102020
rect 442994 102008 443000 102020
rect 443052 102008 443058 102060
rect 147674 100648 147680 100700
rect 147732 100688 147738 100700
rect 256786 100688 256792 100700
rect 147732 100660 256792 100688
rect 147732 100648 147738 100660
rect 256786 100648 256792 100660
rect 256844 100648 256850 100700
rect 342254 100648 342260 100700
rect 342312 100688 342318 100700
rect 438854 100688 438860 100700
rect 342312 100660 438860 100688
rect 342312 100648 342318 100660
rect 438854 100648 438860 100660
rect 438912 100648 438918 100700
rect 150434 100580 150440 100632
rect 150492 100620 150498 100632
rect 256694 100620 256700 100632
rect 150492 100592 256700 100620
rect 150492 100580 150498 100592
rect 256694 100580 256700 100592
rect 256752 100580 256758 100632
rect 342346 100580 342352 100632
rect 342404 100620 342410 100632
rect 434714 100620 434720 100632
rect 342404 100592 434720 100620
rect 342404 100580 342410 100592
rect 434714 100580 434720 100592
rect 434772 100580 434778 100632
rect 145006 99288 145012 99340
rect 145064 99328 145070 99340
rect 256694 99328 256700 99340
rect 145064 99300 256700 99328
rect 145064 99288 145070 99300
rect 256694 99288 256700 99300
rect 256752 99288 256758 99340
rect 342254 99288 342260 99340
rect 342312 99328 342318 99340
rect 430574 99328 430580 99340
rect 342312 99300 430580 99328
rect 342312 99288 342318 99300
rect 430574 99288 430580 99300
rect 430632 99288 430638 99340
rect 138106 97928 138112 97980
rect 138164 97968 138170 97980
rect 256786 97968 256792 97980
rect 138164 97940 256792 97968
rect 138164 97928 138170 97940
rect 256786 97928 256792 97940
rect 256844 97928 256850 97980
rect 342254 97928 342260 97980
rect 342312 97968 342318 97980
rect 425054 97968 425060 97980
rect 342312 97940 425060 97968
rect 342312 97928 342318 97940
rect 425054 97928 425060 97940
rect 425112 97928 425118 97980
rect 140866 97860 140872 97912
rect 140924 97900 140930 97912
rect 256694 97900 256700 97912
rect 140924 97872 256700 97900
rect 140924 97860 140930 97872
rect 256694 97860 256700 97872
rect 256752 97860 256758 97912
rect 342346 97860 342352 97912
rect 342404 97900 342410 97912
rect 420914 97900 420920 97912
rect 342404 97872 420920 97900
rect 342404 97860 342410 97872
rect 420914 97860 420920 97872
rect 420972 97860 420978 97912
rect 132494 96568 132500 96620
rect 132552 96608 132558 96620
rect 256786 96608 256792 96620
rect 132552 96580 256792 96608
rect 132552 96568 132558 96580
rect 256786 96568 256792 96580
rect 256844 96568 256850 96620
rect 342254 96568 342260 96620
rect 342312 96608 342318 96620
rect 416774 96608 416780 96620
rect 342312 96580 416780 96608
rect 342312 96568 342318 96580
rect 416774 96568 416780 96580
rect 416832 96568 416838 96620
rect 135254 96500 135260 96552
rect 135312 96540 135318 96552
rect 256694 96540 256700 96552
rect 135312 96512 256700 96540
rect 135312 96500 135318 96512
rect 256694 96500 256700 96512
rect 256752 96500 256758 96552
rect 342346 96500 342352 96552
rect 342404 96540 342410 96552
rect 412634 96540 412640 96552
rect 342404 96512 412640 96540
rect 342404 96500 342410 96512
rect 412634 96500 412640 96512
rect 412692 96500 412698 96552
rect 129826 95140 129832 95192
rect 129884 95180 129890 95192
rect 256694 95180 256700 95192
rect 129884 95152 256700 95180
rect 129884 95140 129890 95152
rect 256694 95140 256700 95152
rect 256752 95140 256758 95192
rect 342254 95140 342260 95192
rect 342312 95180 342318 95192
rect 395338 95180 395344 95192
rect 342312 95152 395344 95180
rect 342312 95140 342318 95152
rect 395338 95140 395344 95152
rect 395396 95140 395402 95192
rect 122834 93780 122840 93832
rect 122892 93820 122898 93832
rect 256786 93820 256792 93832
rect 122892 93792 256792 93820
rect 122892 93780 122898 93792
rect 256786 93780 256792 93792
rect 256844 93780 256850 93832
rect 342254 93780 342260 93832
rect 342312 93820 342318 93832
rect 402974 93820 402980 93832
rect 342312 93792 402980 93820
rect 342312 93780 342318 93792
rect 402974 93780 402980 93792
rect 403032 93780 403038 93832
rect 125686 93712 125692 93764
rect 125744 93752 125750 93764
rect 256694 93752 256700 93764
rect 125744 93724 256700 93752
rect 125744 93712 125750 93724
rect 256694 93712 256700 93724
rect 256752 93712 256758 93764
rect 342346 93712 342352 93764
rect 342404 93752 342410 93764
rect 398834 93752 398840 93764
rect 342404 93724 398840 93752
rect 342404 93712 342410 93724
rect 398834 93712 398840 93724
rect 398892 93712 398898 93764
rect 117406 92420 117412 92472
rect 117464 92460 117470 92472
rect 256786 92460 256792 92472
rect 117464 92432 256792 92460
rect 117464 92420 117470 92432
rect 256786 92420 256792 92432
rect 256844 92420 256850 92472
rect 342254 92420 342260 92472
rect 342312 92460 342318 92472
rect 394694 92460 394700 92472
rect 342312 92432 394700 92460
rect 342312 92420 342318 92432
rect 394694 92420 394700 92432
rect 394752 92420 394758 92472
rect 120074 92352 120080 92404
rect 120132 92392 120138 92404
rect 256694 92392 256700 92404
rect 120132 92364 256700 92392
rect 120132 92352 120138 92364
rect 256694 92352 256700 92364
rect 256752 92352 256758 92404
rect 342346 92352 342352 92404
rect 342404 92392 342410 92404
rect 389910 92392 389916 92404
rect 342404 92364 389916 92392
rect 342404 92352 342410 92364
rect 389910 92352 389916 92364
rect 389968 92352 389974 92404
rect 209774 90992 209780 91044
rect 209832 91032 209838 91044
rect 256786 91032 256792 91044
rect 209832 91004 256792 91032
rect 209832 90992 209838 91004
rect 256786 90992 256792 91004
rect 256844 90992 256850 91044
rect 342254 90992 342260 91044
rect 342312 91032 342318 91044
rect 522298 91032 522304 91044
rect 342312 91004 522304 91032
rect 342312 90992 342318 91004
rect 522298 90992 522304 91004
rect 522356 90992 522362 91044
rect 212534 90924 212540 90976
rect 212592 90964 212598 90976
rect 256694 90964 256700 90976
rect 212592 90936 256700 90964
rect 212592 90924 212598 90936
rect 256694 90924 256700 90936
rect 256752 90924 256758 90976
rect 342346 90924 342352 90976
rect 342404 90964 342410 90976
rect 520918 90964 520924 90976
rect 342404 90936 520924 90964
rect 342404 90924 342410 90936
rect 520918 90924 520924 90936
rect 520976 90924 520982 90976
rect 207014 89632 207020 89684
rect 207072 89672 207078 89684
rect 256694 89672 256700 89684
rect 207072 89644 256700 89672
rect 207072 89632 207078 89644
rect 256694 89632 256700 89644
rect 256752 89632 256758 89684
rect 342254 89632 342260 89684
rect 342312 89672 342318 89684
rect 519538 89672 519544 89684
rect 342312 89644 519544 89672
rect 342312 89632 342318 89644
rect 519538 89632 519544 89644
rect 519596 89632 519602 89684
rect 200114 88272 200120 88324
rect 200172 88312 200178 88324
rect 256786 88312 256792 88324
rect 200172 88284 256792 88312
rect 200172 88272 200178 88284
rect 256786 88272 256792 88284
rect 256844 88272 256850 88324
rect 342254 88272 342260 88324
rect 342312 88312 342318 88324
rect 514754 88312 514760 88324
rect 342312 88284 514760 88312
rect 342312 88272 342318 88284
rect 514754 88272 514760 88284
rect 514812 88272 514818 88324
rect 204346 88204 204352 88256
rect 204404 88244 204410 88256
rect 256694 88244 256700 88256
rect 204404 88216 256700 88244
rect 204404 88204 204410 88216
rect 256694 88204 256700 88216
rect 256752 88204 256758 88256
rect 342346 88204 342352 88256
rect 342404 88244 342410 88256
rect 510614 88244 510620 88256
rect 342404 88216 510620 88244
rect 342404 88204 342410 88216
rect 510614 88204 510620 88216
rect 510672 88204 510678 88256
rect 194594 86912 194600 86964
rect 194652 86952 194658 86964
rect 256786 86952 256792 86964
rect 194652 86924 256792 86952
rect 194652 86912 194658 86924
rect 256786 86912 256792 86924
rect 256844 86912 256850 86964
rect 342254 86912 342260 86964
rect 342312 86952 342318 86964
rect 506474 86952 506480 86964
rect 342312 86924 506480 86952
rect 342312 86912 342318 86924
rect 506474 86912 506480 86924
rect 506532 86912 506538 86964
rect 197354 86844 197360 86896
rect 197412 86884 197418 86896
rect 256694 86884 256700 86896
rect 197412 86856 256700 86884
rect 197412 86844 197418 86856
rect 256694 86844 256700 86856
rect 256752 86844 256758 86896
rect 342346 86844 342352 86896
rect 342404 86884 342410 86896
rect 502334 86884 502340 86896
rect 342404 86856 502340 86884
rect 342404 86844 342410 86856
rect 502334 86844 502340 86856
rect 502392 86844 502398 86896
rect 187694 85484 187700 85536
rect 187752 85524 187758 85536
rect 256786 85524 256792 85536
rect 187752 85496 256792 85524
rect 187752 85484 187758 85496
rect 256786 85484 256792 85496
rect 256844 85484 256850 85536
rect 342346 85484 342352 85536
rect 342404 85524 342410 85536
rect 492674 85524 492680 85536
rect 342404 85496 492680 85524
rect 342404 85484 342410 85496
rect 492674 85484 492680 85496
rect 492732 85484 492738 85536
rect 191926 85416 191932 85468
rect 191984 85456 191990 85468
rect 256694 85456 256700 85468
rect 191984 85428 256700 85456
rect 191984 85416 191990 85428
rect 256694 85416 256700 85428
rect 256752 85416 256758 85468
rect 342254 85416 342260 85468
rect 342312 85456 342318 85468
rect 465718 85456 465724 85468
rect 342312 85428 465724 85456
rect 342312 85416 342318 85428
rect 465718 85416 465724 85428
rect 465776 85416 465782 85468
rect 184934 84124 184940 84176
rect 184992 84164 184998 84176
rect 256694 84164 256700 84176
rect 184992 84136 256700 84164
rect 184992 84124 184998 84136
rect 256694 84124 256700 84136
rect 256752 84124 256758 84176
rect 342254 84124 342260 84176
rect 342312 84164 342318 84176
rect 488534 84164 488540 84176
rect 342312 84136 488540 84164
rect 342312 84124 342318 84136
rect 488534 84124 488540 84136
rect 488592 84124 488598 84176
rect 179414 82764 179420 82816
rect 179472 82804 179478 82816
rect 256786 82804 256792 82816
rect 179472 82776 256792 82804
rect 179472 82764 179478 82776
rect 256786 82764 256792 82776
rect 256844 82764 256850 82816
rect 342254 82764 342260 82816
rect 342312 82804 342318 82816
rect 484394 82804 484400 82816
rect 342312 82776 484400 82804
rect 342312 82764 342318 82776
rect 484394 82764 484400 82776
rect 484452 82764 484458 82816
rect 182174 82696 182180 82748
rect 182232 82736 182238 82748
rect 256694 82736 256700 82748
rect 182232 82708 256700 82736
rect 182232 82696 182238 82708
rect 256694 82696 256700 82708
rect 256752 82696 256758 82748
rect 342346 82696 342352 82748
rect 342404 82736 342410 82748
rect 461578 82736 461584 82748
rect 342404 82708 461584 82736
rect 342404 82696 342410 82708
rect 461578 82696 461584 82708
rect 461636 82696 461642 82748
rect 172514 81336 172520 81388
rect 172572 81376 172578 81388
rect 256786 81376 256792 81388
rect 172572 81348 256792 81376
rect 172572 81336 172578 81348
rect 256786 81336 256792 81348
rect 256844 81336 256850 81388
rect 342254 81336 342260 81388
rect 342312 81376 342318 81388
rect 476114 81376 476120 81388
rect 342312 81348 476120 81376
rect 342312 81336 342318 81348
rect 476114 81336 476120 81348
rect 476172 81336 476178 81388
rect 176746 81268 176752 81320
rect 176804 81308 176810 81320
rect 256694 81308 256700 81320
rect 176804 81280 256700 81308
rect 176804 81268 176810 81280
rect 256694 81268 256700 81280
rect 256752 81268 256758 81320
rect 342346 81268 342352 81320
rect 342404 81308 342410 81320
rect 470594 81308 470600 81320
rect 342404 81280 470600 81308
rect 342404 81268 342410 81280
rect 470594 81268 470600 81280
rect 470652 81268 470658 81320
rect 166994 79976 167000 80028
rect 167052 80016 167058 80028
rect 256786 80016 256792 80028
rect 167052 79988 256792 80016
rect 167052 79976 167058 79988
rect 256786 79976 256792 79988
rect 256844 79976 256850 80028
rect 342254 79976 342260 80028
rect 342312 80016 342318 80028
rect 466454 80016 466460 80028
rect 342312 79988 466460 80016
rect 342312 79976 342318 79988
rect 466454 79976 466460 79988
rect 466512 79976 466518 80028
rect 169754 79908 169760 79960
rect 169812 79948 169818 79960
rect 256694 79948 256700 79960
rect 169812 79920 256700 79948
rect 169812 79908 169818 79920
rect 256694 79908 256700 79920
rect 256752 79908 256758 79960
rect 342346 79908 342352 79960
rect 342404 79948 342410 79960
rect 453298 79948 453304 79960
rect 342404 79920 453304 79948
rect 342404 79908 342410 79920
rect 453298 79908 453304 79920
rect 453356 79908 453362 79960
rect 164326 78616 164332 78668
rect 164384 78656 164390 78668
rect 256694 78656 256700 78668
rect 164384 78628 256700 78656
rect 164384 78616 164390 78628
rect 256694 78616 256700 78628
rect 256752 78616 256758 78668
rect 342254 78616 342260 78668
rect 342312 78656 342318 78668
rect 458174 78656 458180 78668
rect 342312 78628 458180 78656
rect 342312 78616 342318 78628
rect 458174 78616 458180 78628
rect 458232 78616 458238 78668
rect 157334 77188 157340 77240
rect 157392 77228 157398 77240
rect 256786 77228 256792 77240
rect 157392 77200 256792 77228
rect 157392 77188 157398 77200
rect 256786 77188 256792 77200
rect 256844 77188 256850 77240
rect 342254 77188 342260 77240
rect 342312 77228 342318 77240
rect 454034 77228 454040 77240
rect 342312 77200 454040 77228
rect 342312 77188 342318 77200
rect 454034 77188 454040 77200
rect 454092 77188 454098 77240
rect 161566 77120 161572 77172
rect 161624 77160 161630 77172
rect 256694 77160 256700 77172
rect 161624 77132 256700 77160
rect 161624 77120 161630 77132
rect 256694 77120 256700 77132
rect 256752 77120 256758 77172
rect 342346 77120 342352 77172
rect 342404 77160 342410 77172
rect 448514 77160 448520 77172
rect 342404 77132 448520 77160
rect 342404 77120 342410 77132
rect 448514 77120 448520 77132
rect 448572 77120 448578 77172
rect 151814 75828 151820 75880
rect 151872 75868 151878 75880
rect 256786 75868 256792 75880
rect 151872 75840 256792 75868
rect 151872 75828 151878 75840
rect 256786 75828 256792 75840
rect 256844 75828 256850 75880
rect 342254 75828 342260 75880
rect 342312 75868 342318 75880
rect 443638 75868 443644 75880
rect 342312 75840 443644 75868
rect 342312 75828 342318 75840
rect 443638 75828 443644 75840
rect 443696 75828 443702 75880
rect 154574 75760 154580 75812
rect 154632 75800 154638 75812
rect 256694 75800 256700 75812
rect 154632 75772 256700 75800
rect 154632 75760 154638 75772
rect 256694 75760 256700 75772
rect 256752 75760 256758 75812
rect 342346 75760 342352 75812
rect 342404 75800 342410 75812
rect 440234 75800 440240 75812
rect 342404 75772 440240 75800
rect 342404 75760 342410 75772
rect 440234 75760 440240 75772
rect 440292 75760 440298 75812
rect 149146 74468 149152 74520
rect 149204 74508 149210 74520
rect 256694 74508 256700 74520
rect 149204 74480 256700 74508
rect 149204 74468 149210 74480
rect 256694 74468 256700 74480
rect 256752 74468 256758 74520
rect 342254 74468 342260 74520
rect 342312 74508 342318 74520
rect 436094 74508 436100 74520
rect 342312 74480 436100 74508
rect 342312 74468 342318 74480
rect 436094 74468 436100 74480
rect 436152 74468 436158 74520
rect 142154 73108 142160 73160
rect 142212 73148 142218 73160
rect 256786 73148 256792 73160
rect 142212 73120 256792 73148
rect 142212 73108 142218 73120
rect 256786 73108 256792 73120
rect 256844 73108 256850 73160
rect 342254 73108 342260 73160
rect 342312 73148 342318 73160
rect 431954 73148 431960 73160
rect 342312 73120 431960 73148
rect 342312 73108 342318 73120
rect 431954 73108 431960 73120
rect 432012 73108 432018 73160
rect 144914 73040 144920 73092
rect 144972 73080 144978 73092
rect 256694 73080 256700 73092
rect 144972 73052 256700 73080
rect 144972 73040 144978 73052
rect 256694 73040 256700 73052
rect 256752 73040 256758 73092
rect 342346 73040 342352 73092
rect 342404 73080 342410 73092
rect 417418 73080 417424 73092
rect 342404 73052 417424 73080
rect 342404 73040 342410 73052
rect 417418 73040 417424 73052
rect 417476 73040 417482 73092
rect 136634 71680 136640 71732
rect 136692 71720 136698 71732
rect 256786 71720 256792 71732
rect 136692 71692 256792 71720
rect 136692 71680 136698 71692
rect 256786 71680 256792 71692
rect 256844 71680 256850 71732
rect 342346 71680 342352 71732
rect 342404 71720 342410 71732
rect 418154 71720 418160 71732
rect 342404 71692 418160 71720
rect 342404 71680 342410 71692
rect 418154 71680 418160 71692
rect 418212 71680 418218 71732
rect 139394 71612 139400 71664
rect 139452 71652 139458 71664
rect 256694 71652 256700 71664
rect 139452 71624 256700 71652
rect 139452 71612 139458 71624
rect 256694 71612 256700 71624
rect 256752 71612 256758 71664
rect 342254 71612 342260 71664
rect 342312 71652 342318 71664
rect 413278 71652 413284 71664
rect 342312 71624 413284 71652
rect 342312 71612 342318 71624
rect 413278 71612 413284 71624
rect 413336 71612 413342 71664
rect 129734 70320 129740 70372
rect 129792 70360 129798 70372
rect 256786 70360 256792 70372
rect 129792 70332 256792 70360
rect 129792 70320 129798 70332
rect 256786 70320 256792 70332
rect 256844 70320 256850 70372
rect 342254 70320 342260 70372
rect 342312 70360 342318 70372
rect 414014 70360 414020 70372
rect 342312 70332 414020 70360
rect 342312 70320 342318 70332
rect 414014 70320 414020 70332
rect 414072 70320 414078 70372
rect 133966 70252 133972 70304
rect 134024 70292 134030 70304
rect 256694 70292 256700 70304
rect 134024 70264 256700 70292
rect 134024 70252 134030 70264
rect 256694 70252 256700 70264
rect 256752 70252 256758 70304
rect 342346 70252 342352 70304
rect 342404 70292 342410 70304
rect 409874 70292 409880 70304
rect 342404 70264 409880 70292
rect 342404 70252 342410 70264
rect 409874 70252 409880 70264
rect 409932 70252 409938 70304
rect 126974 68960 126980 69012
rect 127032 69000 127038 69012
rect 256694 69000 256700 69012
rect 127032 68972 256700 69000
rect 127032 68960 127038 68972
rect 256694 68960 256700 68972
rect 256752 68960 256758 69012
rect 342254 68960 342260 69012
rect 342312 69000 342318 69012
rect 399478 69000 399484 69012
rect 342312 68972 399484 69000
rect 342312 68960 342318 68972
rect 399478 68960 399484 68972
rect 399536 68960 399542 69012
rect 121546 67532 121552 67584
rect 121604 67572 121610 67584
rect 256786 67572 256792 67584
rect 121604 67544 256792 67572
rect 121604 67532 121610 67544
rect 256786 67532 256792 67544
rect 256844 67532 256850 67584
rect 342254 67532 342260 67584
rect 342312 67572 342318 67584
rect 400214 67572 400220 67584
rect 342312 67544 400220 67572
rect 342312 67532 342318 67544
rect 400214 67532 400220 67544
rect 400272 67532 400278 67584
rect 124214 67464 124220 67516
rect 124272 67504 124278 67516
rect 256694 67504 256700 67516
rect 124272 67476 256700 67504
rect 124272 67464 124278 67476
rect 256694 67464 256700 67476
rect 256752 67464 256758 67516
rect 342346 67464 342352 67516
rect 342404 67504 342410 67516
rect 396074 67504 396080 67516
rect 342404 67476 396080 67504
rect 342404 67464 342410 67476
rect 396074 67464 396080 67476
rect 396132 67464 396138 67516
rect 117314 66172 117320 66224
rect 117372 66212 117378 66224
rect 256694 66212 256700 66224
rect 117372 66184 256700 66212
rect 117372 66172 117378 66184
rect 256694 66172 256700 66184
rect 256752 66172 256758 66224
rect 342346 66172 342352 66224
rect 342404 66212 342410 66224
rect 482278 66212 482284 66224
rect 342404 66184 482284 66212
rect 342404 66172 342410 66184
rect 482278 66172 482284 66184
rect 482336 66172 482342 66224
rect 211154 66104 211160 66156
rect 211212 66144 211218 66156
rect 256786 66144 256792 66156
rect 211212 66116 256792 66144
rect 211212 66104 211218 66116
rect 256786 66104 256792 66116
rect 256844 66104 256850 66156
rect 342254 66104 342260 66156
rect 342312 66144 342318 66156
rect 391934 66144 391940 66156
rect 342312 66116 391940 66144
rect 342312 66104 342318 66116
rect 391934 66104 391940 66116
rect 391992 66104 391998 66156
rect 208394 64812 208400 64864
rect 208452 64852 208458 64864
rect 256694 64852 256700 64864
rect 208452 64824 256700 64852
rect 208452 64812 208458 64824
rect 256694 64812 256700 64824
rect 256752 64812 256758 64864
rect 342254 64812 342260 64864
rect 342312 64852 342318 64864
rect 475378 64852 475384 64864
rect 342312 64824 475384 64852
rect 342312 64812 342318 64824
rect 475378 64812 475384 64824
rect 475436 64812 475442 64864
rect 201494 63452 201500 63504
rect 201552 63492 201558 63504
rect 256786 63492 256792 63504
rect 201552 63464 256792 63492
rect 201552 63452 201558 63464
rect 256786 63452 256792 63464
rect 256844 63452 256850 63504
rect 342254 63452 342260 63504
rect 342312 63492 342318 63504
rect 472618 63492 472624 63504
rect 342312 63464 472624 63492
rect 342312 63452 342318 63464
rect 472618 63452 472624 63464
rect 472676 63452 472682 63504
rect 204254 63384 204260 63436
rect 204312 63424 204318 63436
rect 256694 63424 256700 63436
rect 204312 63396 256700 63424
rect 204312 63384 204318 63396
rect 256694 63384 256700 63396
rect 256752 63384 256758 63436
rect 342346 63384 342352 63436
rect 342404 63424 342410 63436
rect 468478 63424 468484 63436
rect 342404 63396 468484 63424
rect 342404 63384 342410 63396
rect 468478 63384 468484 63396
rect 468536 63384 468542 63436
rect 195974 62024 195980 62076
rect 196032 62064 196038 62076
rect 256786 62064 256792 62076
rect 196032 62036 256792 62064
rect 196032 62024 196038 62036
rect 256786 62024 256792 62036
rect 256844 62024 256850 62076
rect 342254 62024 342260 62076
rect 342312 62064 342318 62076
rect 464338 62064 464344 62076
rect 342312 62036 464344 62064
rect 342312 62024 342318 62036
rect 464338 62024 464344 62036
rect 464396 62024 464402 62076
rect 198734 61956 198740 62008
rect 198792 61996 198798 62008
rect 256694 61996 256700 62008
rect 198792 61968 256700 61996
rect 198792 61956 198798 61968
rect 256694 61956 256700 61968
rect 256752 61956 256758 62008
rect 342346 61956 342352 62008
rect 342404 61996 342410 62008
rect 460198 61996 460204 62008
rect 342404 61968 460204 61996
rect 342404 61956 342410 61968
rect 460198 61956 460204 61968
rect 460256 61956 460262 62008
rect 189074 60664 189080 60716
rect 189132 60704 189138 60716
rect 256786 60704 256792 60716
rect 189132 60676 256792 60704
rect 189132 60664 189138 60676
rect 256786 60664 256792 60676
rect 256844 60664 256850 60716
rect 342254 60664 342260 60716
rect 342312 60704 342318 60716
rect 450538 60704 450544 60716
rect 342312 60676 450544 60704
rect 342312 60664 342318 60676
rect 450538 60664 450544 60676
rect 450596 60664 450602 60716
rect 191834 60596 191840 60648
rect 191892 60636 191898 60648
rect 256694 60636 256700 60648
rect 191892 60608 256700 60636
rect 191892 60596 191898 60608
rect 256694 60596 256700 60608
rect 256752 60596 256758 60648
rect 342346 60596 342352 60648
rect 342404 60636 342410 60648
rect 446398 60636 446404 60648
rect 342404 60608 446404 60636
rect 342404 60596 342410 60608
rect 446398 60596 446404 60608
rect 446456 60596 446462 60648
rect 186314 59304 186320 59356
rect 186372 59344 186378 59356
rect 256694 59344 256700 59356
rect 186372 59316 256700 59344
rect 186372 59304 186378 59316
rect 256694 59304 256700 59316
rect 256752 59304 256758 59356
rect 342254 59304 342260 59356
rect 342312 59344 342318 59356
rect 489914 59344 489920 59356
rect 342312 59316 489920 59344
rect 342312 59304 342318 59316
rect 489914 59304 489920 59316
rect 489972 59304 489978 59356
rect 180794 57876 180800 57928
rect 180852 57916 180858 57928
rect 256786 57916 256792 57928
rect 180852 57888 256792 57916
rect 180852 57876 180858 57888
rect 256786 57876 256792 57888
rect 256844 57876 256850 57928
rect 342254 57876 342260 57928
rect 342312 57916 342318 57928
rect 485774 57916 485780 57928
rect 342312 57888 485780 57916
rect 342312 57876 342318 57888
rect 485774 57876 485780 57888
rect 485832 57876 485838 57928
rect 183554 57808 183560 57860
rect 183612 57848 183618 57860
rect 256694 57848 256700 57860
rect 183612 57820 256700 57848
rect 183612 57808 183618 57820
rect 256694 57808 256700 57820
rect 256752 57808 256758 57860
rect 342346 57808 342352 57860
rect 342404 57848 342410 57860
rect 481634 57848 481640 57860
rect 342404 57820 481640 57848
rect 342404 57808 342410 57820
rect 481634 57808 481640 57820
rect 481692 57808 481698 57860
rect 173894 56516 173900 56568
rect 173952 56556 173958 56568
rect 256786 56556 256792 56568
rect 173952 56528 256792 56556
rect 173952 56516 173958 56528
rect 256786 56516 256792 56528
rect 256844 56516 256850 56568
rect 342254 56516 342260 56568
rect 342312 56556 342318 56568
rect 477494 56556 477500 56568
rect 342312 56528 477500 56556
rect 342312 56516 342318 56528
rect 477494 56516 477500 56528
rect 477552 56516 477558 56568
rect 176654 56448 176660 56500
rect 176712 56488 176718 56500
rect 256694 56488 256700 56500
rect 176712 56460 256700 56488
rect 176712 56448 176718 56460
rect 256694 56448 256700 56460
rect 256752 56448 256758 56500
rect 342346 56448 342352 56500
rect 342404 56488 342410 56500
rect 471974 56488 471980 56500
rect 342404 56460 471980 56488
rect 342404 56448 342410 56460
rect 471974 56448 471980 56460
rect 472032 56448 472038 56500
rect 171134 55156 171140 55208
rect 171192 55196 171198 55208
rect 256694 55196 256700 55208
rect 171192 55168 256700 55196
rect 171192 55156 171198 55168
rect 256694 55156 256700 55168
rect 256752 55156 256758 55208
rect 342254 55156 342260 55208
rect 342312 55196 342318 55208
rect 467834 55196 467840 55208
rect 342312 55168 467840 55196
rect 342312 55156 342318 55168
rect 467834 55156 467840 55168
rect 467892 55156 467898 55208
rect 164234 53728 164240 53780
rect 164292 53768 164298 53780
rect 256786 53768 256792 53780
rect 164292 53740 256792 53768
rect 164292 53728 164298 53740
rect 256786 53728 256792 53740
rect 256844 53728 256850 53780
rect 342254 53728 342260 53780
rect 342312 53768 342318 53780
rect 463694 53768 463700 53780
rect 342312 53740 463700 53768
rect 342312 53728 342318 53740
rect 463694 53728 463700 53740
rect 463752 53728 463758 53780
rect 168374 53660 168380 53712
rect 168432 53700 168438 53712
rect 256694 53700 256700 53712
rect 168432 53672 256700 53700
rect 168432 53660 168438 53672
rect 256694 53660 256700 53672
rect 256752 53660 256758 53712
rect 342346 53660 342352 53712
rect 342404 53700 342410 53712
rect 459554 53700 459560 53712
rect 342404 53672 459560 53700
rect 342404 53660 342410 53672
rect 459554 53660 459560 53672
rect 459612 53660 459618 53712
rect 158714 52368 158720 52420
rect 158772 52408 158778 52420
rect 256786 52408 256792 52420
rect 158772 52380 256792 52408
rect 158772 52368 158778 52380
rect 256786 52368 256792 52380
rect 256844 52368 256850 52420
rect 342254 52368 342260 52420
rect 342312 52408 342318 52420
rect 455414 52408 455420 52420
rect 342312 52380 455420 52408
rect 342312 52368 342318 52380
rect 455414 52368 455420 52380
rect 455472 52368 455478 52420
rect 161474 52300 161480 52352
rect 161532 52340 161538 52352
rect 256694 52340 256700 52352
rect 161532 52312 256700 52340
rect 161532 52300 161538 52312
rect 256694 52300 256700 52312
rect 256752 52300 256758 52352
rect 342346 52300 342352 52352
rect 342404 52340 342410 52352
rect 449894 52340 449900 52352
rect 342404 52312 449900 52340
rect 342404 52300 342410 52312
rect 449894 52300 449900 52312
rect 449952 52300 449958 52352
rect 153194 51008 153200 51060
rect 153252 51048 153258 51060
rect 256786 51048 256792 51060
rect 153252 51020 256792 51048
rect 153252 51008 153258 51020
rect 256786 51008 256792 51020
rect 256844 51008 256850 51060
rect 342254 51008 342260 51060
rect 342312 51048 342318 51060
rect 445754 51048 445760 51060
rect 342312 51020 445760 51048
rect 342312 51008 342318 51020
rect 445754 51008 445760 51020
rect 445812 51008 445818 51060
rect 155954 50940 155960 50992
rect 156012 50980 156018 50992
rect 256694 50980 256700 50992
rect 156012 50952 256700 50980
rect 156012 50940 156018 50952
rect 256694 50940 256700 50952
rect 256752 50940 256758 50992
rect 342346 50940 342352 50992
rect 342404 50980 342410 50992
rect 441614 50980 441620 50992
rect 342404 50952 441620 50980
rect 342404 50940 342410 50952
rect 441614 50940 441620 50952
rect 441672 50940 441678 50992
rect 149054 49648 149060 49700
rect 149112 49688 149118 49700
rect 256694 49688 256700 49700
rect 149112 49660 256700 49688
rect 149112 49648 149118 49660
rect 256694 49648 256700 49660
rect 256752 49648 256758 49700
rect 342254 49648 342260 49700
rect 342312 49688 342318 49700
rect 437474 49688 437480 49700
rect 342312 49660 437480 49688
rect 342312 49648 342318 49660
rect 437474 49648 437480 49660
rect 437532 49648 437538 49700
rect 143534 48220 143540 48272
rect 143592 48260 143598 48272
rect 256786 48260 256792 48272
rect 143592 48232 256792 48260
rect 143592 48220 143598 48232
rect 256786 48220 256792 48232
rect 256844 48220 256850 48272
rect 342254 48220 342260 48272
rect 342312 48260 342318 48272
rect 433334 48260 433340 48272
rect 342312 48232 433340 48260
rect 342312 48220 342318 48232
rect 433334 48220 433340 48232
rect 433392 48220 433398 48272
rect 146294 48152 146300 48204
rect 146352 48192 146358 48204
rect 256694 48192 256700 48204
rect 146352 48164 256700 48192
rect 146352 48152 146358 48164
rect 256694 48152 256700 48164
rect 256752 48152 256758 48204
rect 342346 48152 342352 48204
rect 342404 48192 342410 48204
rect 427814 48192 427820 48204
rect 342404 48164 427820 48192
rect 342404 48152 342410 48164
rect 427814 48152 427820 48164
rect 427872 48152 427878 48204
rect 138014 46860 138020 46912
rect 138072 46900 138078 46912
rect 256786 46900 256792 46912
rect 138072 46872 256792 46900
rect 138072 46860 138078 46872
rect 256786 46860 256792 46872
rect 256844 46860 256850 46912
rect 342254 46860 342260 46912
rect 342312 46900 342318 46912
rect 423674 46900 423680 46912
rect 342312 46872 423680 46900
rect 342312 46860 342318 46872
rect 423674 46860 423680 46872
rect 423732 46860 423738 46912
rect 140774 46792 140780 46844
rect 140832 46832 140838 46844
rect 256694 46832 256700 46844
rect 140832 46804 256700 46832
rect 140832 46792 140838 46804
rect 256694 46792 256700 46804
rect 256752 46792 256758 46844
rect 342346 46792 342352 46844
rect 342404 46832 342410 46844
rect 358078 46832 358084 46844
rect 342404 46804 358084 46832
rect 342404 46792 342410 46804
rect 358078 46792 358084 46804
rect 358136 46792 358142 46844
rect 131114 45500 131120 45552
rect 131172 45540 131178 45552
rect 256786 45540 256792 45552
rect 131172 45512 256792 45540
rect 131172 45500 131178 45512
rect 256786 45500 256792 45512
rect 256844 45500 256850 45552
rect 342346 45500 342352 45552
rect 342404 45540 342410 45552
rect 411254 45540 411260 45552
rect 342404 45512 411260 45540
rect 342404 45500 342410 45512
rect 411254 45500 411260 45512
rect 411312 45500 411318 45552
rect 133874 45432 133880 45484
rect 133932 45472 133938 45484
rect 256694 45472 256700 45484
rect 133932 45444 256700 45472
rect 133932 45432 133938 45444
rect 256694 45432 256700 45444
rect 256752 45432 256758 45484
rect 342254 45432 342260 45484
rect 342312 45472 342318 45484
rect 388438 45472 388444 45484
rect 342312 45444 388444 45472
rect 342312 45432 342318 45444
rect 388438 45432 388444 45444
rect 388496 45432 388502 45484
rect 128354 44072 128360 44124
rect 128412 44112 128418 44124
rect 256694 44112 256700 44124
rect 128412 44084 256700 44112
rect 128412 44072 128418 44084
rect 256694 44072 256700 44084
rect 256752 44072 256758 44124
rect 342254 44072 342260 44124
rect 342312 44112 342318 44124
rect 405734 44112 405740 44124
rect 342312 44084 405740 44112
rect 342312 44072 342318 44084
rect 405734 44072 405740 44084
rect 405792 44072 405798 44124
rect 121454 42712 121460 42764
rect 121512 42752 121518 42764
rect 256786 42752 256792 42764
rect 121512 42724 256792 42752
rect 121512 42712 121518 42724
rect 256786 42712 256792 42724
rect 256844 42712 256850 42764
rect 342254 42712 342260 42764
rect 342312 42752 342318 42764
rect 382918 42752 382924 42764
rect 342312 42724 382924 42752
rect 342312 42712 342318 42724
rect 382918 42712 382924 42724
rect 382976 42712 382982 42764
rect 125594 42644 125600 42696
rect 125652 42684 125658 42696
rect 256694 42684 256700 42696
rect 125652 42656 256700 42684
rect 125652 42644 125658 42656
rect 256694 42644 256700 42656
rect 256752 42644 256758 42696
rect 342346 42644 342352 42696
rect 342404 42684 342410 42696
rect 381538 42684 381544 42696
rect 342404 42656 381544 42684
rect 342404 42644 342410 42656
rect 381538 42644 381544 42656
rect 381596 42644 381602 42696
rect 115934 41352 115940 41404
rect 115992 41392 115998 41404
rect 256786 41392 256792 41404
rect 115992 41364 256792 41392
rect 115992 41352 115998 41364
rect 256786 41352 256792 41364
rect 256844 41352 256850 41404
rect 342254 41352 342260 41404
rect 342312 41392 342318 41404
rect 389818 41392 389824 41404
rect 342312 41364 389824 41392
rect 342312 41352 342318 41364
rect 389818 41352 389824 41364
rect 389876 41352 389882 41404
rect 118694 41284 118700 41336
rect 118752 41324 118758 41336
rect 256694 41324 256700 41336
rect 118752 41296 256700 41324
rect 118752 41284 118758 41296
rect 256694 41284 256700 41296
rect 256752 41284 256758 41336
rect 342346 41284 342352 41336
rect 342404 41324 342410 41336
rect 389174 41324 389180 41336
rect 342404 41296 389180 41324
rect 342404 41284 342410 41296
rect 389174 41284 389180 41296
rect 389232 41284 389238 41336
rect 124214 38360 124220 38412
rect 124272 38400 124278 38412
rect 336366 38400 336372 38412
rect 124272 38372 336372 38400
rect 124272 38360 124278 38372
rect 336366 38360 336372 38372
rect 336424 38360 336430 38412
rect 106274 38292 106280 38344
rect 106332 38332 106338 38344
rect 332410 38332 332416 38344
rect 106332 38304 332416 38332
rect 106332 38292 106338 38304
rect 332410 38292 332416 38304
rect 332468 38292 332474 38344
rect 99374 38224 99380 38276
rect 99432 38264 99438 38276
rect 330754 38264 330760 38276
rect 99432 38236 330760 38264
rect 99432 38224 99438 38236
rect 330754 38224 330760 38236
rect 330812 38224 330818 38276
rect 50338 38156 50344 38208
rect 50396 38196 50402 38208
rect 316402 38196 316408 38208
rect 50396 38168 316408 38196
rect 50396 38156 50402 38168
rect 316402 38156 316408 38168
rect 316460 38156 316466 38208
rect 51718 38088 51724 38140
rect 51776 38128 51782 38140
rect 317966 38128 317972 38140
rect 51776 38100 317972 38128
rect 51776 38088 51782 38100
rect 317966 38088 317972 38100
rect 318024 38088 318030 38140
rect 35158 38020 35164 38072
rect 35216 38060 35222 38072
rect 314746 38060 314752 38072
rect 35216 38032 314752 38060
rect 35216 38020 35222 38032
rect 314746 38020 314752 38032
rect 314804 38020 314810 38072
rect 320818 38020 320824 38072
rect 320876 38060 320882 38072
rect 320876 38032 321784 38060
rect 320876 38020 320882 38032
rect 22738 37952 22744 38004
rect 22796 37992 22802 38004
rect 313182 37992 313188 38004
rect 22796 37964 313188 37992
rect 22796 37952 22802 37964
rect 313182 37952 313188 37964
rect 313240 37952 313246 38004
rect 318794 37952 318800 38004
rect 318852 37992 318858 38004
rect 319254 37992 319260 38004
rect 318852 37964 319260 37992
rect 318852 37952 318858 37964
rect 319254 37952 319260 37964
rect 319312 37952 319318 38004
rect 320174 37952 320180 38004
rect 320232 37992 320238 38004
rect 320910 37992 320916 38004
rect 320232 37964 320916 37992
rect 320232 37952 320238 37964
rect 320910 37952 320916 37964
rect 320968 37952 320974 38004
rect 321756 37992 321784 38032
rect 322198 38020 322204 38072
rect 322256 38060 322262 38072
rect 337194 38060 337200 38072
rect 322256 38032 337200 38060
rect 322256 38020 322262 38032
rect 337194 38020 337200 38032
rect 337252 38020 337258 38072
rect 334802 37992 334808 38004
rect 321756 37964 334808 37992
rect 334802 37952 334808 37964
rect 334860 37952 334866 38004
rect 10318 37884 10324 37936
rect 10376 37924 10382 37936
rect 337930 37924 337936 37936
rect 10376 37896 318794 37924
rect 10376 37884 10382 37896
rect 264974 37816 264980 37868
rect 265032 37856 265038 37868
rect 265526 37856 265532 37868
rect 265032 37828 265532 37856
rect 265032 37816 265038 37828
rect 265526 37816 265532 37828
rect 265584 37816 265590 37868
rect 266354 37816 266360 37868
rect 266412 37856 266418 37868
rect 267182 37856 267188 37868
rect 266412 37828 267188 37856
rect 266412 37816 266418 37828
rect 267182 37816 267188 37828
rect 267240 37816 267246 37868
rect 270494 37816 270500 37868
rect 270552 37856 270558 37868
rect 271230 37856 271236 37868
rect 270552 37828 271236 37856
rect 270552 37816 270558 37828
rect 271230 37816 271236 37828
rect 271288 37816 271294 37868
rect 274634 37816 274640 37868
rect 274692 37856 274698 37868
rect 275278 37856 275284 37868
rect 274692 37828 275284 37856
rect 274692 37816 274698 37828
rect 275278 37816 275284 37828
rect 275336 37816 275342 37868
rect 276014 37816 276020 37868
rect 276072 37856 276078 37868
rect 276750 37856 276756 37868
rect 276072 37828 276756 37856
rect 276072 37816 276078 37828
rect 276750 37816 276756 37828
rect 276808 37816 276814 37868
rect 318766 37856 318794 37896
rect 328426 37896 337936 37924
rect 328426 37856 328454 37896
rect 337930 37884 337936 37896
rect 337988 37884 337994 37936
rect 318766 37828 328454 37856
rect 271874 36388 271880 36440
rect 271932 36428 271938 36440
rect 272886 36428 272892 36440
rect 271932 36400 272892 36428
rect 271932 36388 271938 36400
rect 272886 36388 272892 36400
rect 272944 36388 272950 36440
rect 321554 35844 321560 35896
rect 321612 35884 321618 35896
rect 322382 35884 322388 35896
rect 321612 35856 322388 35884
rect 321612 35844 321618 35856
rect 322382 35844 322388 35856
rect 322440 35844 322446 35896
rect 120074 21632 120080 21684
rect 120132 21672 120138 21684
rect 335446 21672 335452 21684
rect 120132 21644 335452 21672
rect 120132 21632 120138 21644
rect 335446 21632 335452 21644
rect 335504 21632 335510 21684
rect 113266 21564 113272 21616
rect 113324 21604 113330 21616
rect 334066 21604 334072 21616
rect 113324 21576 334072 21604
rect 113324 21564 113330 21576
rect 334066 21564 334072 21576
rect 334124 21564 334130 21616
rect 110506 21496 110512 21548
rect 110564 21536 110570 21548
rect 332594 21536 332600 21548
rect 110564 21508 332600 21536
rect 110564 21496 110570 21508
rect 332594 21496 332600 21508
rect 332652 21496 332658 21548
rect 102134 21428 102140 21480
rect 102192 21468 102198 21480
rect 331306 21468 331312 21480
rect 102192 21440 331312 21468
rect 102192 21428 102198 21440
rect 331306 21428 331312 21440
rect 331364 21428 331370 21480
rect 45554 21360 45560 21412
rect 45612 21400 45618 21412
rect 318886 21400 318892 21412
rect 45612 21372 318892 21400
rect 45612 21360 45618 21372
rect 318886 21360 318892 21372
rect 318944 21360 318950 21412
rect 95234 20272 95240 20324
rect 95292 20312 95298 20324
rect 329926 20312 329932 20324
rect 95292 20284 329932 20312
rect 95292 20272 95298 20284
rect 329926 20272 329932 20284
rect 329984 20272 329990 20324
rect 92474 20204 92480 20256
rect 92532 20244 92538 20256
rect 328454 20244 328460 20256
rect 92532 20216 328460 20244
rect 92532 20204 92538 20216
rect 328454 20204 328460 20216
rect 328512 20204 328518 20256
rect 88334 20136 88340 20188
rect 88392 20176 88398 20188
rect 327166 20176 327172 20188
rect 88392 20148 327172 20176
rect 88392 20136 88398 20148
rect 327166 20136 327172 20148
rect 327224 20136 327230 20188
rect 85574 20068 85580 20120
rect 85632 20108 85638 20120
rect 327074 20108 327080 20120
rect 85632 20080 327080 20108
rect 85632 20068 85638 20080
rect 327074 20068 327080 20080
rect 327132 20068 327138 20120
rect 81434 20000 81440 20052
rect 81492 20040 81498 20052
rect 325786 20040 325792 20052
rect 81492 20012 325792 20040
rect 81492 20000 81498 20012
rect 325786 20000 325792 20012
rect 325844 20000 325850 20052
rect 13814 19932 13820 19984
rect 13872 19972 13878 19984
rect 311986 19972 311992 19984
rect 13872 19944 311992 19972
rect 13872 19932 13878 19944
rect 311986 19932 311992 19944
rect 312044 19932 312050 19984
rect 77294 18912 77300 18964
rect 77352 18952 77358 18964
rect 325694 18952 325700 18964
rect 77352 18924 325700 18952
rect 77352 18912 77358 18924
rect 325694 18912 325700 18924
rect 325752 18912 325758 18964
rect 74534 18844 74540 18896
rect 74592 18884 74598 18896
rect 324406 18884 324412 18896
rect 74592 18856 324412 18884
rect 74592 18844 74598 18856
rect 324406 18844 324412 18856
rect 324464 18844 324470 18896
rect 70394 18776 70400 18828
rect 70452 18816 70458 18828
rect 324314 18816 324320 18828
rect 70452 18788 324320 18816
rect 70452 18776 70458 18788
rect 324314 18776 324320 18788
rect 324372 18776 324378 18828
rect 67634 18708 67640 18760
rect 67692 18748 67698 18760
rect 322934 18748 322940 18760
rect 67692 18720 322940 18748
rect 67692 18708 67698 18720
rect 322934 18708 322940 18720
rect 322992 18708 322998 18760
rect 63494 18640 63500 18692
rect 63552 18680 63558 18692
rect 321554 18680 321560 18692
rect 63552 18652 321560 18680
rect 63552 18640 63558 18652
rect 321554 18640 321560 18652
rect 321612 18640 321618 18692
rect 60734 18572 60740 18624
rect 60792 18612 60798 18624
rect 321646 18612 321652 18624
rect 60792 18584 321652 18612
rect 60792 18572 60798 18584
rect 321646 18572 321652 18584
rect 321704 18572 321710 18624
rect 44174 17552 44180 17604
rect 44232 17592 44238 17604
rect 292574 17592 292580 17604
rect 44232 17564 292580 17592
rect 44232 17552 44238 17564
rect 292574 17552 292580 17564
rect 292632 17552 292638 17604
rect 41414 17484 41420 17536
rect 41472 17524 41478 17536
rect 291286 17524 291292 17536
rect 41472 17496 291292 17524
rect 41472 17484 41478 17496
rect 291286 17484 291292 17496
rect 291344 17484 291350 17536
rect 56594 17416 56600 17468
rect 56652 17456 56658 17468
rect 320174 17456 320180 17468
rect 56652 17428 320180 17456
rect 56652 17416 56658 17428
rect 320174 17416 320180 17428
rect 320232 17416 320238 17468
rect 52454 17348 52460 17400
rect 52512 17388 52518 17400
rect 320266 17388 320272 17400
rect 52512 17360 320272 17388
rect 52512 17348 52518 17360
rect 320266 17348 320272 17360
rect 320324 17348 320330 17400
rect 49694 17280 49700 17332
rect 49752 17320 49758 17332
rect 318794 17320 318800 17332
rect 49752 17292 318800 17320
rect 49752 17280 49758 17292
rect 318794 17280 318800 17292
rect 318852 17280 318858 17332
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 310606 17252 310612 17264
rect 9732 17224 310612 17252
rect 9732 17212 9738 17224
rect 310606 17212 310612 17224
rect 310664 17212 310670 17264
rect 123018 16260 123024 16312
rect 123076 16300 123082 16312
rect 310514 16300 310520 16312
rect 123076 16272 310520 16300
rect 123076 16260 123082 16272
rect 310514 16260 310520 16272
rect 310572 16260 310578 16312
rect 84194 16192 84200 16244
rect 84252 16232 84258 16244
rect 300946 16232 300952 16244
rect 84252 16204 300952 16232
rect 84252 16192 84258 16204
rect 300946 16192 300952 16204
rect 301004 16192 301010 16244
rect 38378 16124 38384 16176
rect 38436 16164 38442 16176
rect 291194 16164 291200 16176
rect 38436 16136 291200 16164
rect 38436 16124 38442 16136
rect 291194 16124 291200 16136
rect 291252 16124 291258 16176
rect 34514 16056 34520 16108
rect 34572 16096 34578 16108
rect 289906 16096 289912 16108
rect 34572 16068 289912 16096
rect 34572 16056 34578 16068
rect 289906 16056 289912 16068
rect 289964 16056 289970 16108
rect 30834 15988 30840 16040
rect 30892 16028 30898 16040
rect 289814 16028 289820 16040
rect 30892 16000 289820 16028
rect 30892 15988 30898 16000
rect 289814 15988 289820 16000
rect 289872 15988 289878 16040
rect 27706 15920 27712 15972
rect 27764 15960 27770 15972
rect 288434 15960 288440 15972
rect 27764 15932 288440 15960
rect 27764 15920 27770 15932
rect 288434 15920 288440 15932
rect 288492 15920 288498 15972
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 287146 15892 287152 15904
rect 22612 15864 287152 15892
rect 22612 15852 22618 15864
rect 287146 15852 287152 15864
rect 287204 15852 287210 15904
rect 80882 14764 80888 14816
rect 80940 14804 80946 14816
rect 300854 14804 300860 14816
rect 80940 14776 300860 14804
rect 80940 14764 80946 14776
rect 300854 14764 300860 14776
rect 300912 14764 300918 14816
rect 77386 14696 77392 14748
rect 77444 14736 77450 14748
rect 299566 14736 299572 14748
rect 77444 14708 299572 14736
rect 77444 14696 77450 14708
rect 299566 14696 299572 14708
rect 299624 14696 299630 14748
rect 73338 14628 73344 14680
rect 73396 14668 73402 14680
rect 299474 14668 299480 14680
rect 73396 14640 299480 14668
rect 73396 14628 73402 14640
rect 299474 14628 299480 14640
rect 299532 14628 299538 14680
rect 69014 14560 69020 14612
rect 69072 14600 69078 14612
rect 298094 14600 298100 14612
rect 69072 14572 298100 14600
rect 69072 14560 69078 14572
rect 298094 14560 298100 14572
rect 298152 14560 298158 14612
rect 66714 14492 66720 14544
rect 66772 14532 66778 14544
rect 296806 14532 296812 14544
rect 66772 14504 296812 14532
rect 66772 14492 66778 14504
rect 296806 14492 296812 14504
rect 296864 14492 296870 14544
rect 63218 14424 63224 14476
rect 63276 14464 63282 14476
rect 296714 14464 296720 14476
rect 63276 14436 296720 14464
rect 63276 14424 63282 14436
rect 296714 14424 296720 14436
rect 296772 14424 296778 14476
rect 122282 13472 122288 13524
rect 122340 13512 122346 13524
rect 284386 13512 284392 13524
rect 122340 13484 284392 13512
rect 122340 13472 122346 13484
rect 284386 13472 284392 13484
rect 284444 13472 284450 13524
rect 118786 13404 118792 13456
rect 118844 13444 118850 13456
rect 284294 13444 284300 13456
rect 118844 13416 284300 13444
rect 118844 13404 118850 13416
rect 284294 13404 284300 13416
rect 284352 13404 284358 13456
rect 36722 13336 36728 13388
rect 36780 13376 36786 13388
rect 264974 13376 264980 13388
rect 36780 13348 264980 13376
rect 36780 13336 36786 13348
rect 264974 13336 264980 13348
rect 265032 13336 265038 13388
rect 33594 13268 33600 13320
rect 33652 13308 33658 13320
rect 265066 13308 265072 13320
rect 33652 13280 265072 13308
rect 33652 13268 33658 13280
rect 265066 13268 265072 13280
rect 265124 13268 265130 13320
rect 59354 13200 59360 13252
rect 59412 13240 59418 13252
rect 295426 13240 295432 13252
rect 59412 13212 295432 13240
rect 59412 13200 59418 13212
rect 295426 13200 295432 13212
rect 295484 13200 295490 13252
rect 26234 13132 26240 13184
rect 26292 13172 26298 13184
rect 262306 13172 262312 13184
rect 26292 13144 262312 13172
rect 26292 13132 26298 13144
rect 262306 13132 262312 13144
rect 262364 13132 262370 13184
rect 13538 13064 13544 13116
rect 13596 13104 13602 13116
rect 285766 13104 285772 13116
rect 13596 13076 285772 13104
rect 13596 13064 13602 13076
rect 285766 13064 285772 13076
rect 285824 13064 285830 13116
rect 114738 12112 114744 12164
rect 114796 12152 114802 12164
rect 282914 12152 282920 12164
rect 114796 12124 282920 12152
rect 114796 12112 114802 12124
rect 282914 12112 282920 12124
rect 282972 12112 282978 12164
rect 111610 12044 111616 12096
rect 111668 12084 111674 12096
rect 281626 12084 281632 12096
rect 111668 12056 281632 12084
rect 111668 12044 111674 12056
rect 281626 12044 281632 12056
rect 281684 12044 281690 12096
rect 104066 11976 104072 12028
rect 104124 12016 104130 12028
rect 280246 12016 280252 12028
rect 104124 11988 280252 12016
rect 104124 11976 104130 11988
rect 280246 11976 280252 11988
rect 280304 11976 280310 12028
rect 97442 11908 97448 11960
rect 97500 11948 97506 11960
rect 278866 11948 278872 11960
rect 97500 11920 278872 11948
rect 97500 11908 97506 11920
rect 278866 11908 278872 11920
rect 278924 11908 278930 11960
rect 93946 11840 93952 11892
rect 94004 11880 94010 11892
rect 278774 11880 278780 11892
rect 94004 11852 278780 11880
rect 94004 11840 94010 11852
rect 278774 11840 278780 11852
rect 278832 11840 278838 11892
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 262214 11812 262220 11824
rect 21876 11784 262220 11812
rect 21876 11772 21882 11784
rect 262214 11772 262220 11784
rect 262272 11772 262278 11824
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 260926 11744 260932 11756
rect 17092 11716 260932 11744
rect 17092 11704 17098 11716
rect 260926 11704 260932 11716
rect 260984 11704 260990 11756
rect 69106 10616 69112 10668
rect 69164 10656 69170 10668
rect 271874 10656 271880 10668
rect 69164 10628 271880 10656
rect 69164 10616 69170 10628
rect 271874 10616 271880 10628
rect 271932 10616 271938 10668
rect 65058 10548 65064 10600
rect 65116 10588 65122 10600
rect 271966 10588 271972 10600
rect 65116 10560 271972 10588
rect 65116 10548 65122 10560
rect 271966 10548 271972 10560
rect 272024 10548 272030 10600
rect 61562 10480 61568 10532
rect 61620 10520 61626 10532
rect 270494 10520 270500 10532
rect 61620 10492 270500 10520
rect 61620 10480 61626 10492
rect 270494 10480 270500 10492
rect 270552 10480 270558 10532
rect 58434 10412 58440 10464
rect 58492 10452 58498 10464
rect 270586 10452 270592 10464
rect 58492 10424 270592 10452
rect 58492 10412 58498 10424
rect 270586 10412 270592 10424
rect 270644 10412 270650 10464
rect 54938 10344 54944 10396
rect 54996 10384 55002 10396
rect 269206 10384 269212 10396
rect 54996 10356 269212 10384
rect 54996 10344 55002 10356
rect 269206 10344 269212 10356
rect 269264 10344 269270 10396
rect 11882 10276 11888 10328
rect 11940 10316 11946 10328
rect 260834 10316 260840 10328
rect 11940 10288 260840 10316
rect 11940 10276 11946 10288
rect 260834 10276 260840 10288
rect 260892 10276 260898 10328
rect 566 9324 572 9376
rect 624 9364 630 9376
rect 110414 9364 110420 9376
rect 624 9336 110420 9364
rect 624 9324 630 9336
rect 110414 9324 110420 9336
rect 110472 9324 110478 9376
rect 108114 9256 108120 9308
rect 108172 9296 108178 9308
rect 281534 9296 281540 9308
rect 108172 9268 281540 9296
rect 108172 9256 108178 9268
rect 281534 9256 281540 9268
rect 281592 9256 281598 9308
rect 1670 9188 1676 9240
rect 1728 9228 1734 9240
rect 113174 9228 113180 9240
rect 1728 9200 113180 9228
rect 1728 9188 1734 9200
rect 113174 9188 113180 9200
rect 113232 9188 113238 9240
rect 119890 9188 119896 9240
rect 119948 9228 119954 9240
rect 309226 9228 309232 9240
rect 119948 9200 309232 9228
rect 119948 9188 119954 9200
rect 309226 9188 309232 9200
rect 309284 9188 309290 9240
rect 51350 9120 51356 9172
rect 51408 9160 51414 9172
rect 269114 9160 269120 9172
rect 51408 9132 269120 9160
rect 51408 9120 51414 9132
rect 269114 9120 269120 9132
rect 269172 9120 269178 9172
rect 47854 9052 47860 9104
rect 47912 9092 47918 9104
rect 267734 9092 267740 9104
rect 47912 9064 267740 9092
rect 47912 9052 47918 9064
rect 267734 9052 267740 9064
rect 267792 9052 267798 9104
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 259454 9024 259460 9036
rect 7708 8996 259460 9024
rect 7708 8984 7714 8996
rect 259454 8984 259460 8996
rect 259512 8984 259518 9036
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 338114 8956 338120 8968
rect 2924 8928 338120 8956
rect 2924 8916 2930 8928
rect 338114 8916 338120 8928
rect 338172 8916 338178 8968
rect 116394 8168 116400 8220
rect 116452 8208 116458 8220
rect 309134 8208 309140 8220
rect 116452 8180 309140 8208
rect 116452 8168 116458 8180
rect 309134 8168 309140 8180
rect 309192 8168 309198 8220
rect 112806 8100 112812 8152
rect 112864 8140 112870 8152
rect 307754 8140 307760 8152
rect 112864 8112 307760 8140
rect 112864 8100 112870 8112
rect 307754 8100 307760 8112
rect 307812 8100 307818 8152
rect 109310 8032 109316 8084
rect 109368 8072 109374 8084
rect 306466 8072 306472 8084
rect 109368 8044 306472 8072
rect 109368 8032 109374 8044
rect 306466 8032 306472 8044
rect 306524 8032 306530 8084
rect 105722 7964 105728 8016
rect 105780 8004 105786 8016
rect 306374 8004 306380 8016
rect 105780 7976 306380 8004
rect 105780 7964 105786 7976
rect 306374 7964 306380 7976
rect 306432 7964 306438 8016
rect 102226 7896 102232 7948
rect 102284 7936 102290 7948
rect 305086 7936 305092 7948
rect 102284 7908 305092 7936
rect 102284 7896 102290 7908
rect 305086 7896 305092 7908
rect 305144 7896 305150 7948
rect 98638 7828 98644 7880
rect 98696 7868 98702 7880
rect 304994 7868 305000 7880
rect 98696 7840 305000 7868
rect 98696 7828 98702 7840
rect 304994 7828 305000 7840
rect 305052 7828 305058 7880
rect 95142 7760 95148 7812
rect 95200 7800 95206 7812
rect 303614 7800 303620 7812
rect 95200 7772 303620 7800
rect 95200 7760 95206 7772
rect 303614 7760 303620 7772
rect 303672 7760 303678 7812
rect 91554 7692 91560 7744
rect 91612 7732 91618 7744
rect 302326 7732 302332 7744
rect 91612 7704 302332 7732
rect 91612 7692 91618 7704
rect 302326 7692 302332 7704
rect 302384 7692 302390 7744
rect 87966 7624 87972 7676
rect 88024 7664 88030 7676
rect 302234 7664 302240 7676
rect 88024 7636 302240 7664
rect 88024 7624 88030 7636
rect 302234 7624 302240 7636
rect 302292 7624 302298 7676
rect 18230 7556 18236 7608
rect 18288 7596 18294 7608
rect 287054 7596 287060 7608
rect 18288 7568 287060 7596
rect 18288 7556 18294 7568
rect 287054 7556 287060 7568
rect 287112 7556 287118 7608
rect 44266 6604 44272 6656
rect 44324 6644 44330 6656
rect 266354 6644 266360 6656
rect 44324 6616 266360 6644
rect 44324 6604 44330 6616
rect 266354 6604 266360 6616
rect 266412 6604 266418 6656
rect 40678 6536 40684 6588
rect 40736 6576 40742 6588
rect 266446 6576 266452 6588
rect 40736 6548 266452 6576
rect 40736 6536 40742 6548
rect 266446 6536 266452 6548
rect 266504 6536 266510 6588
rect 30098 6468 30104 6520
rect 30156 6508 30162 6520
rect 263594 6508 263600 6520
rect 30156 6480 263600 6508
rect 30156 6468 30162 6480
rect 263594 6468 263600 6480
rect 263652 6468 263658 6520
rect 56042 6400 56048 6452
rect 56100 6440 56106 6452
rect 295334 6440 295340 6452
rect 56100 6412 295340 6440
rect 56100 6400 56106 6412
rect 295334 6400 295340 6412
rect 295392 6400 295398 6452
rect 52546 6332 52552 6384
rect 52604 6372 52610 6384
rect 294046 6372 294052 6384
rect 52604 6344 294052 6372
rect 52604 6332 52610 6344
rect 294046 6332 294052 6344
rect 294104 6332 294110 6384
rect 48958 6264 48964 6316
rect 49016 6304 49022 6316
rect 293954 6304 293960 6316
rect 49016 6276 293960 6304
rect 49016 6264 49022 6276
rect 293954 6264 293960 6276
rect 294012 6264 294018 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 285674 6236 285680 6248
rect 8812 6208 285680 6236
rect 8812 6196 8818 6208
rect 285674 6196 285680 6208
rect 285732 6196 285738 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 339494 6168 339500 6180
rect 4120 6140 339500 6168
rect 4120 6128 4126 6140
rect 339494 6128 339500 6140
rect 339552 6128 339558 6180
rect 101030 5176 101036 5228
rect 101088 5216 101094 5228
rect 280154 5216 280160 5228
rect 101088 5188 280160 5216
rect 101088 5176 101094 5188
rect 280154 5176 280160 5188
rect 280212 5176 280218 5228
rect 90358 5108 90364 5160
rect 90416 5148 90422 5160
rect 277394 5148 277400 5160
rect 90416 5120 277400 5148
rect 90416 5108 90422 5120
rect 277394 5108 277400 5120
rect 277452 5108 277458 5160
rect 86862 5040 86868 5092
rect 86920 5080 86926 5092
rect 276014 5080 276020 5092
rect 86920 5052 276020 5080
rect 86920 5040 86926 5052
rect 276014 5040 276020 5052
rect 276072 5040 276078 5092
rect 83274 4972 83280 5024
rect 83332 5012 83338 5024
rect 276106 5012 276112 5024
rect 83332 4984 276112 5012
rect 83332 4972 83338 4984
rect 276106 4972 276112 4984
rect 276164 4972 276170 5024
rect 79686 4904 79692 4956
rect 79744 4944 79750 4956
rect 274634 4944 274640 4956
rect 79744 4916 274640 4944
rect 79744 4904 79750 4916
rect 274634 4904 274640 4916
rect 274692 4904 274698 4956
rect 76190 4836 76196 4888
rect 76248 4876 76254 4888
rect 274726 4876 274732 4888
rect 76248 4848 274732 4876
rect 76248 4836 76254 4848
rect 274726 4836 274732 4848
rect 274784 4836 274790 4888
rect 72602 4768 72608 4820
rect 72660 4808 72666 4820
rect 273254 4808 273260 4820
rect 72660 4780 273260 4808
rect 72660 4768 72666 4780
rect 273254 4768 273260 4780
rect 273312 4768 273318 4820
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 51718 3788 51724 3800
rect 43128 3760 51724 3788
rect 43128 3748 43134 3760
rect 51718 3748 51724 3760
rect 51776 3748 51782 3800
rect 35986 3680 35992 3732
rect 36044 3720 36050 3732
rect 50338 3720 50344 3732
rect 36044 3692 50344 3720
rect 36044 3680 36050 3692
rect 50338 3680 50344 3692
rect 50396 3680 50402 3732
rect 117590 3680 117596 3732
rect 117648 3720 117654 3732
rect 320818 3720 320824 3732
rect 117648 3692 320824 3720
rect 117648 3680 117654 3692
rect 320818 3680 320824 3692
rect 320876 3680 320882 3732
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 316126 3652 316132 3664
rect 39632 3624 316132 3652
rect 39632 3612 39638 3624
rect 316126 3612 316132 3624
rect 316184 3612 316190 3664
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 314746 3584 314752 3596
rect 32456 3556 314752 3584
rect 32456 3544 32462 3556
rect 314746 3544 314752 3556
rect 314804 3544 314810 3596
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 10318 3516 10324 3528
rect 5316 3488 10324 3516
rect 5316 3476 5322 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 313274 3516 313280 3528
rect 24268 3488 313280 3516
rect 24268 3476 24274 3488
rect 313274 3476 313280 3488
rect 313332 3476 313338 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 322198 3448 322204 3460
rect 6512 3420 322204 3448
rect 6512 3408 6518 3420
rect 322198 3408 322204 3420
rect 322256 3408 322262 3460
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 35158 3380 35164 3392
rect 28960 3352 35164 3380
rect 28960 3340 28966 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 69014 3340 69020 3392
rect 69072 3380 69078 3392
rect 69934 3380 69940 3392
rect 69072 3352 69940 3380
rect 69072 3340 69078 3352
rect 69934 3340 69940 3352
rect 69992 3340 69998 3392
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 22738 3176 22744 3188
rect 19484 3148 22744 3176
rect 19484 3136 19490 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 407120 700408 407172 700460
rect 478512 700408 478564 700460
rect 517520 700408 517572 700460
rect 527180 700408 527232 700460
rect 397460 700340 397512 700392
rect 524420 700340 524472 700392
rect 404360 700272 404412 700324
rect 543464 700272 543516 700324
rect 409880 699660 409932 699712
rect 413652 699660 413704 699712
rect 514760 696940 514812 696992
rect 580172 696940 580224 696992
rect 400220 683136 400272 683188
rect 580172 683136 580224 683188
rect 510620 643084 510672 643136
rect 580172 643084 580224 643136
rect 397460 630640 397512 630692
rect 580172 630640 580224 630692
rect 507860 590656 507912 590708
rect 579804 590656 579856 590708
rect 393320 576852 393372 576904
rect 580172 576852 580224 576904
rect 347780 552712 347832 552764
rect 414020 552712 414072 552764
rect 462320 552712 462372 552764
rect 521660 552712 521712 552764
rect 331220 552644 331272 552696
rect 527916 552644 527968 552696
rect 505744 552440 505796 552492
rect 547144 552440 547196 552492
rect 499212 552372 499264 552424
rect 551284 552372 551336 552424
rect 495992 552304 496044 552356
rect 548524 552304 548576 552356
rect 391664 552236 391716 552288
rect 555424 552236 555476 552288
rect 388352 552168 388404 552220
rect 554044 552168 554096 552220
rect 384948 552100 385000 552152
rect 556804 552100 556856 552152
rect 381912 552032 381964 552084
rect 558184 552032 558236 552084
rect 502340 549244 502392 549296
rect 580264 549244 580316 549296
rect 268384 547884 268436 547936
rect 376944 547884 376996 547936
rect 251824 545096 251876 545148
rect 376944 545096 376996 545148
rect 267004 542376 267056 542428
rect 376852 542376 376904 542428
rect 264244 538228 264296 538280
rect 376944 538228 376996 538280
rect 547144 538160 547196 538212
rect 579896 538160 579948 538212
rect 251916 535440 251968 535492
rect 376944 535440 376996 535492
rect 262864 532720 262916 532772
rect 376944 532720 376996 532772
rect 260104 527144 260156 527196
rect 376944 527144 376996 527196
rect 555424 525716 555476 525768
rect 580172 525716 580224 525768
rect 252008 524424 252060 524476
rect 376944 524424 376996 524476
rect 258724 522996 258776 523048
rect 376944 522996 376996 523048
rect 255964 517488 256016 517540
rect 376944 517488 376996 517540
rect 252100 514768 252152 514820
rect 376944 514768 376996 514820
rect 253204 511980 253256 512032
rect 376944 511980 376996 512032
rect 253296 509260 253348 509312
rect 376944 509260 376996 509312
rect 252468 499468 252520 499520
rect 268384 499468 268436 499520
rect 252468 498108 252520 498160
rect 267004 498108 267056 498160
rect 252468 496748 252520 496800
rect 377404 496748 377456 496800
rect 252376 496680 252428 496732
rect 264244 496680 264296 496732
rect 377312 494708 377364 494760
rect 377772 494708 377824 494760
rect 252376 493960 252428 494012
rect 377496 493960 377548 494012
rect 252468 493892 252520 493944
rect 262864 493892 262916 493944
rect 252468 491988 252520 492040
rect 260104 491988 260156 492040
rect 251824 491308 251876 491360
rect 376944 491308 376996 491360
rect 251916 491172 251968 491224
rect 258724 491172 258776 491224
rect 252468 489812 252520 489864
rect 377588 489812 377640 489864
rect 252008 488520 252060 488572
rect 376944 488520 376996 488572
rect 252468 488452 252520 488504
rect 255964 488452 256016 488504
rect 251916 487160 251968 487212
rect 376944 487160 376996 487212
rect 251272 487092 251324 487144
rect 253204 487092 253256 487144
rect 251732 485732 251784 485784
rect 377680 485732 377732 485784
rect 251364 485596 251416 485648
rect 253296 485596 253348 485648
rect 251732 484304 251784 484356
rect 377312 484304 377364 484356
rect 252468 482944 252520 482996
rect 377864 482944 377916 482996
rect 252376 482876 252428 482928
rect 377956 482876 378008 482928
rect 251732 481584 251784 481636
rect 378048 481584 378100 481636
rect 252468 480156 252520 480208
rect 377404 480156 377456 480208
rect 251732 477436 251784 477488
rect 377496 477436 377548 477488
rect 251916 476076 251968 476128
rect 376944 476076 376996 476128
rect 252468 476008 252520 476060
rect 377220 476008 377272 476060
rect 252468 474648 252520 474700
rect 377036 474648 377088 474700
rect 251548 473356 251600 473408
rect 376944 473356 376996 473408
rect 554044 471928 554096 471980
rect 580172 471928 580224 471980
rect 252468 471248 252520 471300
rect 376944 471248 376996 471300
rect 252468 470500 252520 470552
rect 376944 470500 376996 470552
rect 252468 467780 252520 467832
rect 376944 467780 376996 467832
rect 252376 464992 252428 465044
rect 376944 464992 376996 465044
rect 251272 463768 251324 463820
rect 253204 463768 253256 463820
rect 251548 462272 251600 462324
rect 376944 462272 376996 462324
rect 252468 459484 252520 459536
rect 376944 459484 376996 459536
rect 143448 458056 143500 458108
rect 218704 458056 218756 458108
rect 142068 457988 142120 458040
rect 218796 457988 218848 458040
rect 152464 457920 152516 457972
rect 239128 457920 239180 457972
rect 155224 457852 155276 457904
rect 249156 457852 249208 457904
rect 140044 457784 140096 457836
rect 244832 457784 244884 457836
rect 134524 457716 134576 457768
rect 241980 457716 242032 457768
rect 90364 457648 90416 457700
rect 216312 457648 216364 457700
rect 86224 457580 86276 457632
rect 213460 457580 213512 457632
rect 79324 457512 79376 457564
rect 207756 457512 207808 457564
rect 218888 457512 218940 457564
rect 240600 457512 240652 457564
rect 80704 457444 80756 457496
rect 210608 457444 210660 457496
rect 220084 457444 220136 457496
rect 243452 457444 243504 457496
rect 252284 456696 252336 456748
rect 376944 456696 376996 456748
rect 253204 455336 253256 455388
rect 376944 455336 376996 455388
rect 252192 452548 252244 452600
rect 376852 452548 376904 452600
rect 252008 449828 252060 449880
rect 376944 449828 376996 449880
rect 252100 447040 252152 447092
rect 376944 447040 376996 447092
rect 251916 444320 251968 444372
rect 376852 444320 376904 444372
rect 251824 441532 251876 441584
rect 376944 441532 376996 441584
rect 465724 438676 465776 438728
rect 498200 438676 498252 438728
rect 461584 438608 461636 438660
rect 480352 438608 480404 438660
rect 482284 438608 482336 438660
rect 525892 438608 525944 438660
rect 395344 438540 395396 438592
rect 408500 438540 408552 438592
rect 468484 438540 468536 438592
rect 512644 438540 512696 438592
rect 381544 438472 381596 438524
rect 397920 438472 397972 438524
rect 453304 438472 453356 438524
rect 462596 438472 462648 438524
rect 464344 438472 464396 438524
rect 508228 438472 508280 438524
rect 382924 438404 382976 438456
rect 402336 438404 402388 438456
rect 413284 438404 413336 438456
rect 422944 438404 422996 438456
rect 460204 438404 460256 438456
rect 503812 438404 503864 438456
rect 504364 438404 504416 438456
rect 514116 438404 514168 438456
rect 388444 438336 388496 438388
rect 415584 438336 415636 438388
rect 417424 438336 417476 438388
rect 427360 438336 427412 438388
rect 446404 438336 446456 438388
rect 494980 438336 495032 438388
rect 508504 438336 508556 438388
rect 518532 438336 518584 438388
rect 358084 438268 358136 438320
rect 420000 438268 420052 438320
rect 450544 438268 450596 438320
rect 499580 438268 499632 438320
rect 501604 438268 501656 438320
rect 509700 438268 509752 438320
rect 512644 438268 512696 438320
rect 523040 438268 523092 438320
rect 392584 438200 392636 438252
rect 469956 438200 470008 438252
rect 472624 438200 472676 438252
rect 517060 438200 517112 438252
rect 518164 438200 518216 438252
rect 527364 438200 527416 438252
rect 393964 438132 394016 438184
rect 474372 438132 474424 438184
rect 475384 438132 475436 438184
rect 521660 438132 521712 438184
rect 389824 437520 389876 437572
rect 393504 437520 393556 437572
rect 497464 437520 497516 437572
rect 500960 437520 501012 437572
rect 520924 437520 520976 437572
rect 524420 437520 524472 437572
rect 389916 437452 389968 437504
rect 390560 437452 390612 437504
rect 399484 437452 399536 437504
rect 405280 437452 405332 437504
rect 443644 437452 443696 437504
rect 445024 437452 445076 437504
rect 486424 437452 486476 437504
rect 487620 437452 487672 437504
rect 490564 437452 490616 437504
rect 492036 437452 492088 437504
rect 494704 437452 494756 437504
rect 496452 437452 496504 437504
rect 500224 437452 500276 437504
rect 505284 437452 505336 437504
rect 519544 437452 519596 437504
rect 520280 437452 520332 437504
rect 522304 437452 522356 437504
rect 528836 437452 528888 437504
rect 551284 431876 551336 431928
rect 579804 431876 579856 431928
rect 558184 419432 558236 419484
rect 580172 419432 580224 419484
rect 143448 396992 143500 397044
rect 247040 396992 247092 397044
rect 142068 396924 142120 396976
rect 245660 396924 245712 396976
rect 126888 396856 126940 396908
rect 237380 396856 237432 396908
rect 124128 396788 124180 396840
rect 236000 396788 236052 396840
rect 121368 396720 121420 396772
rect 234620 396720 234672 396772
rect 118608 395632 118660 395684
rect 233240 395632 233292 395684
rect 117228 395564 117280 395616
rect 231860 395564 231912 395616
rect 114468 395496 114520 395548
rect 230480 395496 230532 395548
rect 111708 395428 111760 395480
rect 229100 395428 229152 395480
rect 108948 395360 109000 395412
rect 227720 395360 227772 395412
rect 106188 395292 106240 395344
rect 226340 395292 226392 395344
rect 157340 394272 157392 394324
rect 270500 394272 270552 394324
rect 104808 394204 104860 394256
rect 223580 394204 223632 394256
rect 102048 394136 102100 394188
rect 222200 394136 222252 394188
rect 99288 394068 99340 394120
rect 220820 394068 220872 394120
rect 96528 394000 96580 394052
rect 219440 394000 219492 394052
rect 93768 393932 93820 393984
rect 218060 393932 218112 393984
rect 149060 392980 149112 393032
rect 255320 392980 255372 393032
rect 150440 392912 150492 392964
rect 258264 392912 258316 392964
rect 151820 392844 151872 392896
rect 260840 392844 260892 392896
rect 153200 392776 153252 392828
rect 263600 392776 263652 392828
rect 154580 392708 154632 392760
rect 264980 392708 265032 392760
rect 155960 392640 156012 392692
rect 268108 392640 268160 392692
rect 71320 392572 71372 392624
rect 205640 392572 205692 392624
rect 147680 391620 147732 391672
rect 252560 391620 252612 391672
rect 158720 391552 158772 391604
rect 273260 391552 273312 391604
rect 161480 391484 161532 391536
rect 277952 391484 278004 391536
rect 160100 391416 160152 391468
rect 276020 391416 276072 391468
rect 162860 391348 162912 391400
rect 280160 391348 280212 391400
rect 68744 391280 68796 391332
rect 204260 391280 204312 391332
rect 189080 391212 189132 391264
rect 325884 391212 325936 391264
rect 159824 390192 159876 390244
rect 191840 390192 191892 390244
rect 158536 390124 158588 390176
rect 193220 390124 193272 390176
rect 144920 390056 144972 390108
rect 248512 390056 248564 390108
rect 186320 389988 186372 390040
rect 320180 389988 320232 390040
rect 132500 389920 132552 389972
rect 338120 389920 338172 389972
rect 131120 389852 131172 389904
rect 339500 389852 339552 389904
rect 129740 389784 129792 389836
rect 359280 389784 359332 389836
rect 176660 388832 176712 388884
rect 305000 388832 305052 388884
rect 178040 388764 178092 388816
rect 307760 388764 307812 388816
rect 179420 388696 179472 388748
rect 310520 388696 310572 388748
rect 180800 388628 180852 388680
rect 313280 388628 313332 388680
rect 183560 388560 183612 388612
rect 317420 388560 317472 388612
rect 182180 388492 182232 388544
rect 316040 388492 316092 388544
rect 187700 388424 187752 388476
rect 322940 388424 322992 388476
rect 146300 387676 146352 387728
rect 249800 387676 249852 387728
rect 164240 387608 164292 387660
rect 282920 387608 282972 387660
rect 165620 387540 165672 387592
rect 285680 387540 285732 387592
rect 167000 387472 167052 387524
rect 288440 387472 288492 387524
rect 168380 387404 168432 387456
rect 289820 387404 289872 387456
rect 169760 387336 169812 387388
rect 292580 387336 292632 387388
rect 171140 387268 171192 387320
rect 295340 387268 295392 387320
rect 172520 387200 172572 387252
rect 298100 387200 298152 387252
rect 175280 387132 175332 387184
rect 302240 387132 302292 387184
rect 173900 387064 173952 387116
rect 300860 387064 300912 387116
rect 78496 386316 78548 386368
rect 80704 386316 80756 386368
rect 89168 386316 89220 386368
rect 90364 386316 90416 386368
rect 133696 386316 133748 386368
rect 134524 386316 134576 386368
rect 138480 386316 138532 386368
rect 140044 386316 140096 386368
rect 146208 386316 146260 386368
rect 155224 386316 155276 386368
rect 73896 386248 73948 386300
rect 79324 386248 79376 386300
rect 81072 386248 81124 386300
rect 211160 386248 211212 386300
rect 86500 386180 86552 386232
rect 213920 386180 213972 386232
rect 92112 386112 92164 386164
rect 216680 386112 216732 386164
rect 131028 386044 131080 386096
rect 218888 386044 218940 386096
rect 136088 385976 136140 386028
rect 220084 385976 220136 386028
rect 128636 385908 128688 385960
rect 152464 385908 152516 385960
rect 77208 385840 77260 385892
rect 208400 385840 208452 385892
rect 351000 385636 351052 385688
rect 380900 385636 380952 385688
rect 83648 385092 83700 385144
rect 86224 385092 86276 385144
rect 170864 384616 170916 384668
rect 177304 384616 177356 384668
rect 217876 384616 217928 384668
rect 351000 384616 351052 384668
rect 139400 384548 139452 384600
rect 358820 384548 358872 384600
rect 138020 384480 138072 384532
rect 358912 384480 358964 384532
rect 136640 384412 136692 384464
rect 359004 384412 359056 384464
rect 135260 384344 135312 384396
rect 359096 384344 359148 384396
rect 133880 384276 133932 384328
rect 359188 384276 359240 384328
rect 178684 379448 178736 379500
rect 190460 379448 190512 379500
rect 548524 379448 548576 379500
rect 580172 379448 580224 379500
rect 556804 365644 556856 365696
rect 580172 365644 580224 365696
rect 176660 336744 176712 336796
rect 216680 336744 216732 336796
rect 178684 320084 178736 320136
rect 194600 320084 194652 320136
rect 178960 318724 179012 318776
rect 195980 318724 196032 318776
rect 178960 317364 179012 317416
rect 197360 317364 197412 317416
rect 178592 315936 178644 315988
rect 198740 315936 198792 315988
rect 178684 314576 178736 314628
rect 200120 314576 200172 314628
rect 182824 309136 182876 309188
rect 216680 309136 216732 309188
rect 177304 309068 177356 309120
rect 216772 309068 216824 309120
rect 39120 299412 39172 299464
rect 39948 299412 40000 299464
rect 177304 299412 177356 299464
rect 163228 298868 163280 298920
rect 201500 298868 201552 298920
rect 163412 298732 163464 298784
rect 202880 298732 202932 298784
rect 218704 298052 218756 298104
rect 343364 298052 343416 298104
rect 136088 297984 136140 298036
rect 140044 297984 140096 298036
rect 218796 297984 218848 298036
rect 343180 297984 343232 298036
rect 264336 297916 264388 297968
rect 265348 297916 265400 297968
rect 275284 297916 275336 297968
rect 276756 297916 276808 297968
rect 282184 297916 282236 297968
rect 285956 297916 286008 297968
rect 287704 297916 287756 297968
rect 295340 297916 295392 297968
rect 68836 297848 68888 297900
rect 69664 297848 69716 297900
rect 77208 297304 77260 297356
rect 259552 297304 259604 297356
rect 203524 297236 203576 297288
rect 238116 297236 238168 297288
rect 108580 297168 108632 297220
rect 125876 297168 125928 297220
rect 141056 297168 141108 297220
rect 162124 297168 162176 297220
rect 202144 297168 202196 297220
rect 276020 297168 276072 297220
rect 108948 297100 109000 297152
rect 251548 297100 251600 297152
rect 108856 297032 108908 297084
rect 259460 297032 259512 297084
rect 302884 297032 302936 297084
rect 315764 297032 315816 297084
rect 108672 296964 108724 297016
rect 269764 296964 269816 297016
rect 294604 296964 294656 297016
rect 302332 296964 302384 297016
rect 305644 296964 305696 297016
rect 320916 296964 320968 297016
rect 86224 296896 86276 296948
rect 259460 296896 259512 296948
rect 289084 296896 289136 296948
rect 298468 296896 298520 296948
rect 300124 296896 300176 296948
rect 310980 296896 311032 296948
rect 83372 296828 83424 296880
rect 259736 296828 259788 296880
rect 295984 296828 296036 296880
rect 305092 296828 305144 296880
rect 80704 296760 80756 296812
rect 259644 296760 259696 296812
rect 286324 296760 286376 296812
rect 290004 296760 290056 296812
rect 291844 296760 291896 296812
rect 300860 296760 300912 296812
rect 304264 296760 304316 296812
rect 317420 296760 317472 296812
rect 108764 296692 108816 296744
rect 117412 296692 117464 296744
rect 129648 296692 129700 296744
rect 137284 296692 137336 296744
rect 264244 296692 264296 296744
rect 268016 296692 268068 296744
rect 284944 296692 284996 296744
rect 287612 296692 287664 296744
rect 298744 296692 298796 296744
rect 308588 296692 308640 296744
rect 205640 296012 205692 296064
rect 261116 296012 261168 296064
rect 198740 295944 198792 295996
rect 260196 295944 260248 295996
rect 160100 242156 160152 242208
rect 260932 242156 260984 242208
rect 191840 240932 191892 240984
rect 280160 240932 280212 240984
rect 109224 240864 109276 240916
rect 292580 240864 292632 240916
rect 73068 240796 73120 240848
rect 260196 240796 260248 240848
rect 109592 240728 109644 240780
rect 313280 240728 313332 240780
rect 71688 239368 71740 239420
rect 260104 239368 260156 239420
rect 89628 238076 89680 238128
rect 229836 238076 229888 238128
rect 90916 238008 90968 238060
rect 233332 238008 233384 238060
rect 174728 236988 174780 237040
rect 251364 236988 251416 237040
rect 167736 236920 167788 236972
rect 249800 236920 249852 236972
rect 157248 236852 157300 236904
rect 248420 236852 248472 236904
rect 82728 236784 82780 236836
rect 208952 236784 209004 236836
rect 244188 236784 244240 236836
rect 273444 236784 273496 236836
rect 84016 236716 84068 236768
rect 222936 236716 222988 236768
rect 240968 236716 241020 236768
rect 271880 236716 271932 236768
rect 77116 236648 77168 236700
rect 260288 236648 260340 236700
rect 38936 235560 38988 235612
rect 111340 235560 111392 235612
rect 188620 235560 188672 235612
rect 258172 235560 258224 235612
rect 79968 235492 80020 235544
rect 194968 235492 195020 235544
rect 216588 235492 216640 235544
rect 262220 235492 262272 235544
rect 109040 235424 109092 235476
rect 255320 235424 255372 235476
rect 109132 235356 109184 235408
rect 256700 235356 256752 235408
rect 109316 235288 109368 235340
rect 265072 235288 265124 235340
rect 109408 235220 109460 235272
rect 267832 235220 267884 235272
rect 57888 234132 57940 234184
rect 132592 234132 132644 234184
rect 136364 234132 136416 234184
rect 217508 234132 217560 234184
rect 38844 234064 38896 234116
rect 139400 234064 139452 234116
rect 170956 234064 171008 234116
rect 217324 234064 217376 234116
rect 39028 233996 39080 234048
rect 146300 233996 146352 234048
rect 150256 233996 150308 234048
rect 247040 233996 247092 234048
rect 56508 233928 56560 233980
rect 118240 233928 118292 233980
rect 129372 233928 129424 233980
rect 236000 233928 236052 233980
rect 38292 233860 38344 233912
rect 181076 233860 181128 233912
rect 77024 233044 77076 233096
rect 142712 233044 142764 233096
rect 115388 232976 115440 233028
rect 182824 232976 182876 233028
rect 185216 232976 185268 233028
rect 202144 232976 202196 233028
rect 125876 232908 125928 232960
rect 203524 232908 203576 232960
rect 213092 232908 213144 232960
rect 284944 232908 284996 232960
rect 81256 232840 81308 232892
rect 163596 232840 163648 232892
rect 202604 232840 202656 232892
rect 282184 232840 282236 232892
rect 68836 232772 68888 232824
rect 153200 232772 153252 232824
rect 162124 232772 162176 232824
rect 258172 232772 258224 232824
rect 137284 232704 137336 232756
rect 236828 232704 236880 232756
rect 242808 232704 242860 232756
rect 261116 232704 261168 232756
rect 68744 232636 68796 232688
rect 121736 232636 121788 232688
rect 140044 232636 140096 232688
rect 247316 232636 247368 232688
rect 251088 232636 251140 232688
rect 260840 232636 260892 232688
rect 111708 232568 111760 232620
rect 219624 232568 219676 232620
rect 254952 232568 255004 232620
rect 275284 232568 275336 232620
rect 114468 232500 114520 232552
rect 226340 232500 226392 232552
rect 251456 232500 251508 232552
rect 304264 232500 304316 232552
rect 217968 231752 218020 231804
rect 262680 231752 262732 231804
rect 139308 231684 139360 231736
rect 262956 231684 263008 231736
rect 133788 231616 133840 231668
rect 262864 231616 262916 231668
rect 124128 231548 124180 231600
rect 262772 231548 262824 231600
rect 109500 231480 109552 231532
rect 115940 231480 115992 231532
rect 121368 231480 121420 231532
rect 261300 231480 261352 231532
rect 108212 231412 108264 231464
rect 252560 231412 252612 231464
rect 256608 231412 256660 231464
rect 261208 231412 261260 231464
rect 108304 231344 108356 231396
rect 258080 231344 258132 231396
rect 91008 231276 91060 231328
rect 262404 231276 262456 231328
rect 108488 231208 108540 231260
rect 322940 231208 322992 231260
rect 60556 231140 60608 231192
rect 261024 231140 261076 231192
rect 110328 231072 110380 231124
rect 325700 231072 325752 231124
rect 237288 231004 237340 231056
rect 260472 231004 260524 231056
rect 240048 230936 240100 230988
rect 260564 230936 260616 230988
rect 146208 230392 146260 230444
rect 259368 230392 259420 230444
rect 217876 230052 217928 230104
rect 263048 230052 263100 230104
rect 248328 229984 248380 230036
rect 260012 229984 260064 230036
rect 99196 229916 99248 229968
rect 259920 229916 259972 229968
rect 108396 229848 108448 229900
rect 262588 229848 262640 229900
rect 99104 229780 99156 229832
rect 259828 229780 259880 229832
rect 96436 229712 96488 229764
rect 262496 229712 262548 229764
rect 263508 224884 263560 224936
rect 276664 224884 276716 224936
rect 261116 224272 261168 224324
rect 259828 224204 259880 224256
rect 260472 224204 260524 224256
rect 262312 224204 262364 224256
rect 262680 224204 262732 224256
rect 261116 224068 261168 224120
rect 262772 223864 262824 223916
rect 262772 223660 262824 223712
rect 97908 223524 97960 223576
rect 107660 223524 107712 223576
rect 262956 223524 263008 223576
rect 305644 223524 305696 223576
rect 260012 222164 260064 222216
rect 260564 222164 260616 222216
rect 93676 217948 93728 218000
rect 107660 217948 107712 218000
rect 263508 217948 263560 218000
rect 300124 217948 300176 218000
rect 263508 216588 263560 216640
rect 298744 216588 298796 216640
rect 263508 213868 263560 213920
rect 294604 213868 294656 213920
rect 263508 211080 263560 211132
rect 291844 211080 291896 211132
rect 263508 204212 263560 204264
rect 277492 204212 277544 204264
rect 262220 189932 262272 189984
rect 264336 189932 264388 189984
rect 75828 188980 75880 189032
rect 107660 188980 107712 189032
rect 88156 186260 88208 186312
rect 107660 186260 107712 186312
rect 38752 180752 38804 180804
rect 107660 180752 107712 180804
rect 78496 177964 78548 178016
rect 107660 177964 107712 178016
rect 62028 172456 62080 172508
rect 107660 172456 107712 172508
rect 74448 169668 74500 169720
rect 107660 169668 107712 169720
rect 63408 164160 63460 164212
rect 107660 164160 107712 164212
rect 38476 161372 38528 161424
rect 107660 161372 107712 161424
rect 96528 160420 96580 160472
rect 110604 160420 110656 160472
rect 260380 160080 260432 160132
rect 263692 160080 263744 160132
rect 242808 159400 242860 159452
rect 273352 159400 273404 159452
rect 110420 159332 110472 159384
rect 111156 159332 111208 159384
rect 244280 159332 244332 159384
rect 282920 159332 282972 159384
rect 85488 159264 85540 159316
rect 240692 159264 240744 159316
rect 78588 159196 78640 159248
rect 233516 159196 233568 159248
rect 256608 159196 256660 159248
rect 274640 159196 274692 159248
rect 86776 159128 86828 159180
rect 243728 159128 243780 159180
rect 246396 159128 246448 159180
rect 266452 159128 266504 159180
rect 92296 159060 92348 159112
rect 249892 159060 249944 159112
rect 253572 159060 253624 159112
rect 273260 159060 273312 159112
rect 95148 158992 95200 159044
rect 253940 158992 253992 159044
rect 259368 158992 259420 159044
rect 278780 158992 278832 159044
rect 88248 158924 88300 158976
rect 247132 158924 247184 158976
rect 249524 158924 249576 158976
rect 270592 158924 270644 158976
rect 38660 158856 38712 158908
rect 217232 158856 217284 158908
rect 243360 158856 243412 158908
rect 266360 158856 266412 158908
rect 38568 158788 38620 158840
rect 224316 158788 224368 158840
rect 240048 158788 240100 158840
rect 263600 158788 263652 158840
rect 39948 158720 40000 158772
rect 110420 158720 110472 158772
rect 113180 158720 113232 158772
rect 383660 158720 383712 158772
rect 60648 158652 60700 158704
rect 219440 158652 219492 158704
rect 235908 158652 235960 158704
rect 244280 158652 244332 158704
rect 248236 158652 248288 158704
rect 295984 158652 296036 158704
rect 92388 158584 92440 158636
rect 251272 158584 251324 158636
rect 255596 158584 255648 158636
rect 302884 158584 302936 158636
rect 69664 158516 69716 158568
rect 225328 158516 225380 158568
rect 239312 158516 239364 158568
rect 286324 158516 286376 158568
rect 59268 158448 59320 158500
rect 214196 158448 214248 158500
rect 242348 158448 242400 158500
rect 287704 158448 287756 158500
rect 67548 158380 67600 158432
rect 221280 158380 221332 158432
rect 231124 158380 231176 158432
rect 242808 158380 242860 158432
rect 245384 158380 245436 158432
rect 289084 158380 289136 158432
rect 110604 158312 110656 158364
rect 256976 158312 257028 158364
rect 230112 158244 230164 158296
rect 270500 158244 270552 158296
rect 227076 158176 227128 158228
rect 260380 158176 260432 158228
rect 102048 158108 102100 158160
rect 234620 158108 234672 158160
rect 104808 158040 104860 158092
rect 236552 158040 236604 158092
rect 106188 157972 106240 158024
rect 237656 157972 237708 158024
rect 228088 157904 228140 157956
rect 264244 157904 264296 157956
rect 99288 157836 99340 157888
rect 232504 157836 232556 157888
rect 93768 157768 93820 157820
rect 231860 157768 231912 157820
rect 114560 155932 114612 155984
rect 115204 155932 115256 155984
rect 117320 155932 117372 155984
rect 118240 155932 118292 155984
rect 121460 155932 121512 155984
rect 122380 155932 122432 155984
rect 129740 155932 129792 155984
rect 130476 155932 130528 155984
rect 133880 155932 133932 155984
rect 134616 155932 134668 155984
rect 144920 155932 144972 155984
rect 145840 155932 145892 155984
rect 149060 155932 149112 155984
rect 149888 155932 149940 155984
rect 157340 155932 157392 155984
rect 158076 155932 158128 155984
rect 161480 155932 161532 155984
rect 162124 155932 162176 155984
rect 164240 155932 164292 155984
rect 165160 155932 165212 155984
rect 172520 155932 172572 155984
rect 173348 155932 173400 155984
rect 176660 155932 176712 155984
rect 177396 155932 177448 155984
rect 184940 155932 184992 155984
rect 185584 155932 185636 155984
rect 187700 155932 187752 155984
rect 188620 155932 188672 155984
rect 200120 155932 200172 155984
rect 200856 155932 200908 155984
rect 204260 155932 204312 155984
rect 204996 155932 205048 155984
rect 191840 153688 191892 153740
rect 192760 153688 192812 153740
rect 111800 120028 111852 120080
rect 256700 120028 256752 120080
rect 342260 120028 342312 120080
rect 382280 120028 382332 120080
rect 110512 118600 110564 118652
rect 256700 118600 256752 118652
rect 342352 118600 342404 118652
rect 386420 118600 386472 118652
rect 114652 118532 114704 118584
rect 256792 118532 256844 118584
rect 342260 118532 342312 118584
rect 379520 118532 379572 118584
rect 114560 117240 114612 117292
rect 256700 117240 256752 117292
rect 342352 117240 342404 117292
rect 518164 117240 518216 117292
rect 211252 117172 211304 117224
rect 256792 117172 256844 117224
rect 342260 117172 342312 117224
rect 387800 117172 387852 117224
rect 205640 115880 205692 115932
rect 256792 115880 256844 115932
rect 342260 115880 342312 115932
rect 512644 115880 512696 115932
rect 208492 115812 208544 115864
rect 256700 115812 256752 115864
rect 342352 115812 342404 115864
rect 508504 115812 508556 115864
rect 202880 114452 202932 114504
rect 256700 114452 256752 114504
rect 342260 114452 342312 114504
rect 504364 114452 504416 114504
rect 196072 113092 196124 113144
rect 256792 113092 256844 113144
rect 342260 113092 342312 113144
rect 501604 113092 501656 113144
rect 200212 113024 200264 113076
rect 256700 113024 256752 113076
rect 342352 113024 342404 113076
rect 500224 113024 500276 113076
rect 190460 111732 190512 111784
rect 256792 111732 256844 111784
rect 342260 111732 342312 111784
rect 497464 111732 497516 111784
rect 193220 111664 193272 111716
rect 256700 111664 256752 111716
rect 342352 111664 342404 111716
rect 494704 111664 494756 111716
rect 187792 110372 187844 110424
rect 256700 110372 256752 110424
rect 342260 110372 342312 110424
rect 490564 110372 490616 110424
rect 180892 108944 180944 108996
rect 256792 108944 256844 108996
rect 342260 108944 342312 108996
rect 486424 108944 486476 108996
rect 185032 108876 185084 108928
rect 256700 108876 256752 108928
rect 342352 108876 342404 108928
rect 483020 108876 483072 108928
rect 175280 107584 175332 107636
rect 256792 107584 256844 107636
rect 342260 107584 342312 107636
rect 478880 107584 478932 107636
rect 178040 107516 178092 107568
rect 256700 107516 256752 107568
rect 342352 107516 342404 107568
rect 393964 107516 394016 107568
rect 168472 106224 168524 106276
rect 256792 106224 256844 106276
rect 342352 106224 342404 106276
rect 465080 106224 465132 106276
rect 172612 106156 172664 106208
rect 256700 106156 256752 106208
rect 342260 106156 342312 106208
rect 392584 106156 392636 106208
rect 165620 104796 165672 104848
rect 256700 104796 256752 104848
rect 342260 104796 342312 104848
rect 460940 104796 460992 104848
rect 160100 103436 160152 103488
rect 256792 103436 256844 103488
rect 342260 103436 342312 103488
rect 456800 103436 456852 103488
rect 162860 103368 162912 103420
rect 256700 103368 256752 103420
rect 342352 103368 342404 103420
rect 452660 103368 452712 103420
rect 153292 102076 153344 102128
rect 256792 102076 256844 102128
rect 342260 102076 342312 102128
rect 447140 102076 447192 102128
rect 157432 102008 157484 102060
rect 256700 102008 256752 102060
rect 342352 102008 342404 102060
rect 443000 102008 443052 102060
rect 147680 100648 147732 100700
rect 256792 100648 256844 100700
rect 342260 100648 342312 100700
rect 438860 100648 438912 100700
rect 150440 100580 150492 100632
rect 256700 100580 256752 100632
rect 342352 100580 342404 100632
rect 434720 100580 434772 100632
rect 145012 99288 145064 99340
rect 256700 99288 256752 99340
rect 342260 99288 342312 99340
rect 430580 99288 430632 99340
rect 138112 97928 138164 97980
rect 256792 97928 256844 97980
rect 342260 97928 342312 97980
rect 425060 97928 425112 97980
rect 140872 97860 140924 97912
rect 256700 97860 256752 97912
rect 342352 97860 342404 97912
rect 420920 97860 420972 97912
rect 132500 96568 132552 96620
rect 256792 96568 256844 96620
rect 342260 96568 342312 96620
rect 416780 96568 416832 96620
rect 135260 96500 135312 96552
rect 256700 96500 256752 96552
rect 342352 96500 342404 96552
rect 412640 96500 412692 96552
rect 129832 95140 129884 95192
rect 256700 95140 256752 95192
rect 342260 95140 342312 95192
rect 395344 95140 395396 95192
rect 122840 93780 122892 93832
rect 256792 93780 256844 93832
rect 342260 93780 342312 93832
rect 402980 93780 403032 93832
rect 125692 93712 125744 93764
rect 256700 93712 256752 93764
rect 342352 93712 342404 93764
rect 398840 93712 398892 93764
rect 117412 92420 117464 92472
rect 256792 92420 256844 92472
rect 342260 92420 342312 92472
rect 394700 92420 394752 92472
rect 120080 92352 120132 92404
rect 256700 92352 256752 92404
rect 342352 92352 342404 92404
rect 389916 92352 389968 92404
rect 209780 90992 209832 91044
rect 256792 90992 256844 91044
rect 342260 90992 342312 91044
rect 522304 90992 522356 91044
rect 212540 90924 212592 90976
rect 256700 90924 256752 90976
rect 342352 90924 342404 90976
rect 520924 90924 520976 90976
rect 207020 89632 207072 89684
rect 256700 89632 256752 89684
rect 342260 89632 342312 89684
rect 519544 89632 519596 89684
rect 200120 88272 200172 88324
rect 256792 88272 256844 88324
rect 342260 88272 342312 88324
rect 514760 88272 514812 88324
rect 204352 88204 204404 88256
rect 256700 88204 256752 88256
rect 342352 88204 342404 88256
rect 510620 88204 510672 88256
rect 194600 86912 194652 86964
rect 256792 86912 256844 86964
rect 342260 86912 342312 86964
rect 506480 86912 506532 86964
rect 197360 86844 197412 86896
rect 256700 86844 256752 86896
rect 342352 86844 342404 86896
rect 502340 86844 502392 86896
rect 187700 85484 187752 85536
rect 256792 85484 256844 85536
rect 342352 85484 342404 85536
rect 492680 85484 492732 85536
rect 191932 85416 191984 85468
rect 256700 85416 256752 85468
rect 342260 85416 342312 85468
rect 465724 85416 465776 85468
rect 184940 84124 184992 84176
rect 256700 84124 256752 84176
rect 342260 84124 342312 84176
rect 488540 84124 488592 84176
rect 179420 82764 179472 82816
rect 256792 82764 256844 82816
rect 342260 82764 342312 82816
rect 484400 82764 484452 82816
rect 182180 82696 182232 82748
rect 256700 82696 256752 82748
rect 342352 82696 342404 82748
rect 461584 82696 461636 82748
rect 172520 81336 172572 81388
rect 256792 81336 256844 81388
rect 342260 81336 342312 81388
rect 476120 81336 476172 81388
rect 176752 81268 176804 81320
rect 256700 81268 256752 81320
rect 342352 81268 342404 81320
rect 470600 81268 470652 81320
rect 167000 79976 167052 80028
rect 256792 79976 256844 80028
rect 342260 79976 342312 80028
rect 466460 79976 466512 80028
rect 169760 79908 169812 79960
rect 256700 79908 256752 79960
rect 342352 79908 342404 79960
rect 453304 79908 453356 79960
rect 164332 78616 164384 78668
rect 256700 78616 256752 78668
rect 342260 78616 342312 78668
rect 458180 78616 458232 78668
rect 157340 77188 157392 77240
rect 256792 77188 256844 77240
rect 342260 77188 342312 77240
rect 454040 77188 454092 77240
rect 161572 77120 161624 77172
rect 256700 77120 256752 77172
rect 342352 77120 342404 77172
rect 448520 77120 448572 77172
rect 151820 75828 151872 75880
rect 256792 75828 256844 75880
rect 342260 75828 342312 75880
rect 443644 75828 443696 75880
rect 154580 75760 154632 75812
rect 256700 75760 256752 75812
rect 342352 75760 342404 75812
rect 440240 75760 440292 75812
rect 149152 74468 149204 74520
rect 256700 74468 256752 74520
rect 342260 74468 342312 74520
rect 436100 74468 436152 74520
rect 142160 73108 142212 73160
rect 256792 73108 256844 73160
rect 342260 73108 342312 73160
rect 431960 73108 432012 73160
rect 144920 73040 144972 73092
rect 256700 73040 256752 73092
rect 342352 73040 342404 73092
rect 417424 73040 417476 73092
rect 136640 71680 136692 71732
rect 256792 71680 256844 71732
rect 342352 71680 342404 71732
rect 418160 71680 418212 71732
rect 139400 71612 139452 71664
rect 256700 71612 256752 71664
rect 342260 71612 342312 71664
rect 413284 71612 413336 71664
rect 129740 70320 129792 70372
rect 256792 70320 256844 70372
rect 342260 70320 342312 70372
rect 414020 70320 414072 70372
rect 133972 70252 134024 70304
rect 256700 70252 256752 70304
rect 342352 70252 342404 70304
rect 409880 70252 409932 70304
rect 126980 68960 127032 69012
rect 256700 68960 256752 69012
rect 342260 68960 342312 69012
rect 399484 68960 399536 69012
rect 121552 67532 121604 67584
rect 256792 67532 256844 67584
rect 342260 67532 342312 67584
rect 400220 67532 400272 67584
rect 124220 67464 124272 67516
rect 256700 67464 256752 67516
rect 342352 67464 342404 67516
rect 396080 67464 396132 67516
rect 117320 66172 117372 66224
rect 256700 66172 256752 66224
rect 342352 66172 342404 66224
rect 482284 66172 482336 66224
rect 211160 66104 211212 66156
rect 256792 66104 256844 66156
rect 342260 66104 342312 66156
rect 391940 66104 391992 66156
rect 208400 64812 208452 64864
rect 256700 64812 256752 64864
rect 342260 64812 342312 64864
rect 475384 64812 475436 64864
rect 201500 63452 201552 63504
rect 256792 63452 256844 63504
rect 342260 63452 342312 63504
rect 472624 63452 472676 63504
rect 204260 63384 204312 63436
rect 256700 63384 256752 63436
rect 342352 63384 342404 63436
rect 468484 63384 468536 63436
rect 195980 62024 196032 62076
rect 256792 62024 256844 62076
rect 342260 62024 342312 62076
rect 464344 62024 464396 62076
rect 198740 61956 198792 62008
rect 256700 61956 256752 62008
rect 342352 61956 342404 62008
rect 460204 61956 460256 62008
rect 189080 60664 189132 60716
rect 256792 60664 256844 60716
rect 342260 60664 342312 60716
rect 450544 60664 450596 60716
rect 191840 60596 191892 60648
rect 256700 60596 256752 60648
rect 342352 60596 342404 60648
rect 446404 60596 446456 60648
rect 186320 59304 186372 59356
rect 256700 59304 256752 59356
rect 342260 59304 342312 59356
rect 489920 59304 489972 59356
rect 180800 57876 180852 57928
rect 256792 57876 256844 57928
rect 342260 57876 342312 57928
rect 485780 57876 485832 57928
rect 183560 57808 183612 57860
rect 256700 57808 256752 57860
rect 342352 57808 342404 57860
rect 481640 57808 481692 57860
rect 173900 56516 173952 56568
rect 256792 56516 256844 56568
rect 342260 56516 342312 56568
rect 477500 56516 477552 56568
rect 176660 56448 176712 56500
rect 256700 56448 256752 56500
rect 342352 56448 342404 56500
rect 471980 56448 472032 56500
rect 171140 55156 171192 55208
rect 256700 55156 256752 55208
rect 342260 55156 342312 55208
rect 467840 55156 467892 55208
rect 164240 53728 164292 53780
rect 256792 53728 256844 53780
rect 342260 53728 342312 53780
rect 463700 53728 463752 53780
rect 168380 53660 168432 53712
rect 256700 53660 256752 53712
rect 342352 53660 342404 53712
rect 459560 53660 459612 53712
rect 158720 52368 158772 52420
rect 256792 52368 256844 52420
rect 342260 52368 342312 52420
rect 455420 52368 455472 52420
rect 161480 52300 161532 52352
rect 256700 52300 256752 52352
rect 342352 52300 342404 52352
rect 449900 52300 449952 52352
rect 153200 51008 153252 51060
rect 256792 51008 256844 51060
rect 342260 51008 342312 51060
rect 445760 51008 445812 51060
rect 155960 50940 156012 50992
rect 256700 50940 256752 50992
rect 342352 50940 342404 50992
rect 441620 50940 441672 50992
rect 149060 49648 149112 49700
rect 256700 49648 256752 49700
rect 342260 49648 342312 49700
rect 437480 49648 437532 49700
rect 143540 48220 143592 48272
rect 256792 48220 256844 48272
rect 342260 48220 342312 48272
rect 433340 48220 433392 48272
rect 146300 48152 146352 48204
rect 256700 48152 256752 48204
rect 342352 48152 342404 48204
rect 427820 48152 427872 48204
rect 138020 46860 138072 46912
rect 256792 46860 256844 46912
rect 342260 46860 342312 46912
rect 423680 46860 423732 46912
rect 140780 46792 140832 46844
rect 256700 46792 256752 46844
rect 342352 46792 342404 46844
rect 358084 46792 358136 46844
rect 131120 45500 131172 45552
rect 256792 45500 256844 45552
rect 342352 45500 342404 45552
rect 411260 45500 411312 45552
rect 133880 45432 133932 45484
rect 256700 45432 256752 45484
rect 342260 45432 342312 45484
rect 388444 45432 388496 45484
rect 128360 44072 128412 44124
rect 256700 44072 256752 44124
rect 342260 44072 342312 44124
rect 405740 44072 405792 44124
rect 121460 42712 121512 42764
rect 256792 42712 256844 42764
rect 342260 42712 342312 42764
rect 382924 42712 382976 42764
rect 125600 42644 125652 42696
rect 256700 42644 256752 42696
rect 342352 42644 342404 42696
rect 381544 42644 381596 42696
rect 115940 41352 115992 41404
rect 256792 41352 256844 41404
rect 342260 41352 342312 41404
rect 389824 41352 389876 41404
rect 118700 41284 118752 41336
rect 256700 41284 256752 41336
rect 342352 41284 342404 41336
rect 389180 41284 389232 41336
rect 124220 38360 124272 38412
rect 336372 38360 336424 38412
rect 106280 38292 106332 38344
rect 332416 38292 332468 38344
rect 99380 38224 99432 38276
rect 330760 38224 330812 38276
rect 50344 38156 50396 38208
rect 316408 38156 316460 38208
rect 51724 38088 51776 38140
rect 317972 38088 318024 38140
rect 35164 38020 35216 38072
rect 314752 38020 314804 38072
rect 320824 38020 320876 38072
rect 22744 37952 22796 38004
rect 313188 37952 313240 38004
rect 318800 37952 318852 38004
rect 319260 37952 319312 38004
rect 320180 37952 320232 38004
rect 320916 37952 320968 38004
rect 322204 38020 322256 38072
rect 337200 38020 337252 38072
rect 334808 37952 334860 38004
rect 10324 37884 10376 37936
rect 264980 37816 265032 37868
rect 265532 37816 265584 37868
rect 266360 37816 266412 37868
rect 267188 37816 267240 37868
rect 270500 37816 270552 37868
rect 271236 37816 271288 37868
rect 274640 37816 274692 37868
rect 275284 37816 275336 37868
rect 276020 37816 276072 37868
rect 276756 37816 276808 37868
rect 337936 37884 337988 37936
rect 271880 36388 271932 36440
rect 272892 36388 272944 36440
rect 321560 35844 321612 35896
rect 322388 35844 322440 35896
rect 120080 21632 120132 21684
rect 335452 21632 335504 21684
rect 113272 21564 113324 21616
rect 334072 21564 334124 21616
rect 110512 21496 110564 21548
rect 332600 21496 332652 21548
rect 102140 21428 102192 21480
rect 331312 21428 331364 21480
rect 45560 21360 45612 21412
rect 318892 21360 318944 21412
rect 95240 20272 95292 20324
rect 329932 20272 329984 20324
rect 92480 20204 92532 20256
rect 328460 20204 328512 20256
rect 88340 20136 88392 20188
rect 327172 20136 327224 20188
rect 85580 20068 85632 20120
rect 327080 20068 327132 20120
rect 81440 20000 81492 20052
rect 325792 20000 325844 20052
rect 13820 19932 13872 19984
rect 311992 19932 312044 19984
rect 77300 18912 77352 18964
rect 325700 18912 325752 18964
rect 74540 18844 74592 18896
rect 324412 18844 324464 18896
rect 70400 18776 70452 18828
rect 324320 18776 324372 18828
rect 67640 18708 67692 18760
rect 322940 18708 322992 18760
rect 63500 18640 63552 18692
rect 321560 18640 321612 18692
rect 60740 18572 60792 18624
rect 321652 18572 321704 18624
rect 44180 17552 44232 17604
rect 292580 17552 292632 17604
rect 41420 17484 41472 17536
rect 291292 17484 291344 17536
rect 56600 17416 56652 17468
rect 320180 17416 320232 17468
rect 52460 17348 52512 17400
rect 320272 17348 320324 17400
rect 49700 17280 49752 17332
rect 318800 17280 318852 17332
rect 9680 17212 9732 17264
rect 310612 17212 310664 17264
rect 123024 16260 123076 16312
rect 310520 16260 310572 16312
rect 84200 16192 84252 16244
rect 300952 16192 301004 16244
rect 38384 16124 38436 16176
rect 291200 16124 291252 16176
rect 34520 16056 34572 16108
rect 289912 16056 289964 16108
rect 30840 15988 30892 16040
rect 289820 15988 289872 16040
rect 27712 15920 27764 15972
rect 288440 15920 288492 15972
rect 22560 15852 22612 15904
rect 287152 15852 287204 15904
rect 80888 14764 80940 14816
rect 300860 14764 300912 14816
rect 77392 14696 77444 14748
rect 299572 14696 299624 14748
rect 73344 14628 73396 14680
rect 299480 14628 299532 14680
rect 69020 14560 69072 14612
rect 298100 14560 298152 14612
rect 66720 14492 66772 14544
rect 296812 14492 296864 14544
rect 63224 14424 63276 14476
rect 296720 14424 296772 14476
rect 122288 13472 122340 13524
rect 284392 13472 284444 13524
rect 118792 13404 118844 13456
rect 284300 13404 284352 13456
rect 36728 13336 36780 13388
rect 264980 13336 265032 13388
rect 33600 13268 33652 13320
rect 265072 13268 265124 13320
rect 59360 13200 59412 13252
rect 295432 13200 295484 13252
rect 26240 13132 26292 13184
rect 262312 13132 262364 13184
rect 13544 13064 13596 13116
rect 285772 13064 285824 13116
rect 114744 12112 114796 12164
rect 282920 12112 282972 12164
rect 111616 12044 111668 12096
rect 281632 12044 281684 12096
rect 104072 11976 104124 12028
rect 280252 11976 280304 12028
rect 97448 11908 97500 11960
rect 278872 11908 278924 11960
rect 93952 11840 94004 11892
rect 278780 11840 278832 11892
rect 21824 11772 21876 11824
rect 262220 11772 262272 11824
rect 17040 11704 17092 11756
rect 260932 11704 260984 11756
rect 69112 10616 69164 10668
rect 271880 10616 271932 10668
rect 65064 10548 65116 10600
rect 271972 10548 272024 10600
rect 61568 10480 61620 10532
rect 270500 10480 270552 10532
rect 58440 10412 58492 10464
rect 270592 10412 270644 10464
rect 54944 10344 54996 10396
rect 269212 10344 269264 10396
rect 11888 10276 11940 10328
rect 260840 10276 260892 10328
rect 572 9324 624 9376
rect 110420 9324 110472 9376
rect 108120 9256 108172 9308
rect 281540 9256 281592 9308
rect 1676 9188 1728 9240
rect 113180 9188 113232 9240
rect 119896 9188 119948 9240
rect 309232 9188 309284 9240
rect 51356 9120 51408 9172
rect 269120 9120 269172 9172
rect 47860 9052 47912 9104
rect 267740 9052 267792 9104
rect 7656 8984 7708 9036
rect 259460 8984 259512 9036
rect 2872 8916 2924 8968
rect 338120 8916 338172 8968
rect 116400 8168 116452 8220
rect 309140 8168 309192 8220
rect 112812 8100 112864 8152
rect 307760 8100 307812 8152
rect 109316 8032 109368 8084
rect 306472 8032 306524 8084
rect 105728 7964 105780 8016
rect 306380 7964 306432 8016
rect 102232 7896 102284 7948
rect 305092 7896 305144 7948
rect 98644 7828 98696 7880
rect 305000 7828 305052 7880
rect 95148 7760 95200 7812
rect 303620 7760 303672 7812
rect 91560 7692 91612 7744
rect 302332 7692 302384 7744
rect 87972 7624 88024 7676
rect 302240 7624 302292 7676
rect 18236 7556 18288 7608
rect 287060 7556 287112 7608
rect 44272 6604 44324 6656
rect 266360 6604 266412 6656
rect 40684 6536 40736 6588
rect 266452 6536 266504 6588
rect 30104 6468 30156 6520
rect 263600 6468 263652 6520
rect 56048 6400 56100 6452
rect 295340 6400 295392 6452
rect 52552 6332 52604 6384
rect 294052 6332 294104 6384
rect 48964 6264 49016 6316
rect 293960 6264 294012 6316
rect 8760 6196 8812 6248
rect 285680 6196 285732 6248
rect 4068 6128 4120 6180
rect 339500 6128 339552 6180
rect 101036 5176 101088 5228
rect 280160 5176 280212 5228
rect 90364 5108 90416 5160
rect 277400 5108 277452 5160
rect 86868 5040 86920 5092
rect 276020 5040 276072 5092
rect 83280 4972 83332 5024
rect 276112 4972 276164 5024
rect 79692 4904 79744 4956
rect 274640 4904 274692 4956
rect 76196 4836 76248 4888
rect 274732 4836 274784 4888
rect 72608 4768 72660 4820
rect 273260 4768 273312 4820
rect 43076 3748 43128 3800
rect 51724 3748 51776 3800
rect 35992 3680 36044 3732
rect 50344 3680 50396 3732
rect 117596 3680 117648 3732
rect 320824 3680 320876 3732
rect 39580 3612 39632 3664
rect 316132 3612 316184 3664
rect 32404 3544 32456 3596
rect 314752 3544 314804 3596
rect 5264 3476 5316 3528
rect 10324 3476 10376 3528
rect 24216 3476 24268 3528
rect 313280 3476 313332 3528
rect 6460 3408 6512 3460
rect 322204 3408 322256 3460
rect 28908 3340 28960 3392
rect 35164 3340 35216 3392
rect 69020 3340 69072 3392
rect 69940 3340 69992 3392
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 19432 3136 19484 3188
rect 22744 3136 22796 3188
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 552702 331260 702986
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 347792 552770 347820 702406
rect 397472 700398 397500 703520
rect 407120 700460 407172 700466
rect 407120 700402 407172 700408
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 404360 700324 404412 700330
rect 404360 700266 404412 700272
rect 400220 683188 400272 683194
rect 400220 683130 400272 683136
rect 397460 630692 397512 630698
rect 397460 630634 397512 630640
rect 393320 576904 393372 576910
rect 393320 576846 393372 576852
rect 393332 557534 393360 576846
rect 393332 557506 394188 557534
rect 347780 552764 347832 552770
rect 347780 552706 347832 552712
rect 331220 552696 331272 552702
rect 331220 552638 331272 552644
rect 391664 552288 391716 552294
rect 391664 552230 391716 552236
rect 388352 552220 388404 552226
rect 388352 552162 388404 552168
rect 384948 552152 385000 552158
rect 384948 552094 385000 552100
rect 381912 552084 381964 552090
rect 381912 552026 381964 552032
rect 381924 549930 381952 552026
rect 384960 549930 384988 552094
rect 388364 549930 388392 552162
rect 391676 549930 391704 552230
rect 381616 549902 381952 549930
rect 384836 549902 384988 549930
rect 388056 549902 388392 549930
rect 391368 549902 391704 549930
rect 394160 549930 394188 557506
rect 397472 549930 397500 630634
rect 400232 557534 400260 683130
rect 400232 557506 400720 557534
rect 400692 549930 400720 557506
rect 404372 549930 404400 700266
rect 407132 557534 407160 700402
rect 413664 699718 413692 703520
rect 409880 699712 409932 699718
rect 409880 699654 409932 699660
rect 413652 699712 413704 699718
rect 413652 699654 413704 699660
rect 409892 557534 409920 699654
rect 407132 557506 407252 557534
rect 409892 557506 410472 557534
rect 407224 549930 407252 557506
rect 410444 549930 410472 557506
rect 462332 552770 462360 703520
rect 478524 700466 478552 703520
rect 527192 700466 527220 703520
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 517520 700460 517572 700466
rect 517520 700402 517572 700408
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 514760 696992 514812 696998
rect 514760 696934 514812 696940
rect 510620 643136 510672 643142
rect 510620 643078 510672 643084
rect 507860 590708 507912 590714
rect 507860 590650 507912 590656
rect 507872 557534 507900 590650
rect 510632 557534 510660 643078
rect 507872 557506 508268 557534
rect 510632 557506 511580 557534
rect 414020 552764 414072 552770
rect 414020 552706 414072 552712
rect 462320 552764 462372 552770
rect 462320 552706 462372 552712
rect 414032 549930 414060 552706
rect 505744 552492 505796 552498
rect 505744 552434 505796 552440
rect 499212 552424 499264 552430
rect 499212 552366 499264 552372
rect 495992 552356 496044 552362
rect 495992 552298 496044 552304
rect 496004 549930 496032 552298
rect 499224 549930 499252 552366
rect 505756 549930 505784 552434
rect 394160 549902 394588 549930
rect 397472 549902 397900 549930
rect 400692 549902 401120 549930
rect 404372 549902 404432 549930
rect 407224 549902 407652 549930
rect 410444 549902 410872 549930
rect 414032 549902 414184 549930
rect 495696 549902 496032 549930
rect 498916 549902 499252 549930
rect 505448 549902 505784 549930
rect 508240 549930 508268 557506
rect 511552 549930 511580 557506
rect 514772 549930 514800 696934
rect 517532 557534 517560 700402
rect 524420 700392 524472 700398
rect 524420 700334 524472 700340
rect 524432 557534 524460 700334
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 517532 557506 518112 557534
rect 524432 557506 524644 557534
rect 518084 549930 518112 557506
rect 521660 552764 521712 552770
rect 521660 552706 521712 552712
rect 521672 549930 521700 552706
rect 524616 549930 524644 557506
rect 527916 552696 527968 552702
rect 527916 552638 527968 552644
rect 527928 549930 527956 552638
rect 547144 552492 547196 552498
rect 547144 552434 547196 552440
rect 508240 549902 508668 549930
rect 511552 549902 511980 549930
rect 514772 549902 515200 549930
rect 518084 549902 518512 549930
rect 521672 549902 521732 549930
rect 524616 549902 525044 549930
rect 527928 549902 528264 549930
rect 502228 549358 502380 549386
rect 502352 549302 502380 549358
rect 502340 549296 502392 549302
rect 502340 549238 502392 549244
rect 376942 548720 376998 548729
rect 376942 548655 376998 548664
rect 376956 547942 376984 548655
rect 268384 547936 268436 547942
rect 268384 547878 268436 547884
rect 376944 547936 376996 547942
rect 376944 547878 376996 547884
rect 251824 545148 251876 545154
rect 251824 545090 251876 545096
rect 251836 499089 251864 545090
rect 267004 542428 267056 542434
rect 267004 542370 267056 542376
rect 264244 538280 264296 538286
rect 264244 538222 264296 538228
rect 251916 535492 251968 535498
rect 251916 535434 251968 535440
rect 251822 499080 251878 499089
rect 251822 499015 251878 499024
rect 251928 495281 251956 535434
rect 262864 532772 262916 532778
rect 262864 532714 262916 532720
rect 260104 527196 260156 527202
rect 260104 527138 260156 527144
rect 252008 524476 252060 524482
rect 252008 524418 252060 524424
rect 251914 495272 251970 495281
rect 251914 495207 251970 495216
rect 251824 491360 251876 491366
rect 251824 491302 251876 491308
rect 251272 487144 251324 487150
rect 251272 487086 251324 487092
rect 251284 486985 251312 487086
rect 251270 486976 251326 486985
rect 251270 486911 251326 486920
rect 251732 485784 251784 485790
rect 251732 485726 251784 485732
rect 251364 485648 251416 485654
rect 251362 485616 251364 485625
rect 251416 485616 251418 485625
rect 251362 485551 251418 485560
rect 251744 485081 251772 485726
rect 251730 485072 251786 485081
rect 251730 485007 251786 485016
rect 251732 484356 251784 484362
rect 251732 484298 251784 484304
rect 251744 483993 251772 484298
rect 251730 483984 251786 483993
rect 251730 483919 251786 483928
rect 251732 481636 251784 481642
rect 251732 481578 251784 481584
rect 251744 481273 251772 481578
rect 251730 481264 251786 481273
rect 251730 481199 251786 481208
rect 251836 479505 251864 491302
rect 251916 491224 251968 491230
rect 252020 491201 252048 524418
rect 258724 523048 258776 523054
rect 258724 522990 258776 522996
rect 255964 517540 256016 517546
rect 255964 517482 256016 517488
rect 252100 514820 252152 514826
rect 252100 514762 252152 514768
rect 251916 491166 251968 491172
rect 252006 491192 252062 491201
rect 251928 490657 251956 491166
rect 252006 491127 252062 491136
rect 251914 490648 251970 490657
rect 251914 490583 251970 490592
rect 252008 488572 252060 488578
rect 252008 488514 252060 488520
rect 251916 487212 251968 487218
rect 251916 487154 251968 487160
rect 251822 479496 251878 479505
rect 251822 479431 251878 479440
rect 251732 477488 251784 477494
rect 251928 477465 251956 487154
rect 252020 478553 252048 488514
rect 252112 487937 252140 514762
rect 253204 512032 253256 512038
rect 253204 511974 253256 511980
rect 252468 499520 252520 499526
rect 252468 499462 252520 499468
rect 252480 499361 252508 499462
rect 252466 499352 252522 499361
rect 252466 499287 252522 499296
rect 252468 498160 252520 498166
rect 252468 498102 252520 498108
rect 252480 497865 252508 498102
rect 252466 497856 252522 497865
rect 252466 497791 252522 497800
rect 252468 496800 252520 496806
rect 252466 496768 252468 496777
rect 252520 496768 252522 496777
rect 252376 496732 252428 496738
rect 252466 496703 252522 496712
rect 252376 496674 252428 496680
rect 252388 496233 252416 496674
rect 252374 496224 252430 496233
rect 252374 496159 252430 496168
rect 252466 494048 252522 494057
rect 252376 494012 252428 494018
rect 252466 493983 252522 493992
rect 252376 493954 252428 493960
rect 252388 493513 252416 493954
rect 252480 493950 252508 493983
rect 252468 493944 252520 493950
rect 252468 493886 252520 493892
rect 252374 493504 252430 493513
rect 252374 493439 252430 493448
rect 252466 492144 252522 492153
rect 252466 492079 252522 492088
rect 252480 492046 252508 492079
rect 252468 492040 252520 492046
rect 252468 491982 252520 491988
rect 252468 489864 252520 489870
rect 252468 489806 252520 489812
rect 252480 489569 252508 489806
rect 252466 489560 252522 489569
rect 252466 489495 252522 489504
rect 252468 488504 252520 488510
rect 252466 488472 252468 488481
rect 252520 488472 252522 488481
rect 252466 488407 252522 488416
rect 252098 487928 252154 487937
rect 252098 487863 252154 487872
rect 253216 487150 253244 511974
rect 253296 509312 253348 509318
rect 253296 509254 253348 509260
rect 253204 487144 253256 487150
rect 253204 487086 253256 487092
rect 253308 485654 253336 509254
rect 255976 488510 256004 517482
rect 258736 491230 258764 522990
rect 260116 492046 260144 527138
rect 262876 493950 262904 532714
rect 264256 496738 264284 538222
rect 267016 498166 267044 542370
rect 268396 499526 268424 547878
rect 376942 546136 376998 546145
rect 376942 546071 376998 546080
rect 376956 545154 376984 546071
rect 376944 545148 376996 545154
rect 376944 545090 376996 545096
rect 376850 543552 376906 543561
rect 376850 543487 376906 543496
rect 376864 542434 376892 543487
rect 376852 542428 376904 542434
rect 376852 542370 376904 542376
rect 377402 540968 377458 540977
rect 377402 540903 377458 540912
rect 376942 538384 376998 538393
rect 376942 538319 376998 538328
rect 376956 538286 376984 538319
rect 376944 538280 376996 538286
rect 376944 538222 376996 538228
rect 376942 535936 376998 535945
rect 376942 535871 376998 535880
rect 376956 535498 376984 535871
rect 376944 535492 376996 535498
rect 376944 535434 376996 535440
rect 376942 533352 376998 533361
rect 376942 533287 376998 533296
rect 376956 532778 376984 533287
rect 376944 532772 376996 532778
rect 376944 532714 376996 532720
rect 376942 528184 376998 528193
rect 376942 528119 376998 528128
rect 376956 527202 376984 528119
rect 376944 527196 376996 527202
rect 376944 527138 376996 527144
rect 376942 525600 376998 525609
rect 376942 525535 376998 525544
rect 376956 524482 376984 525535
rect 376944 524476 376996 524482
rect 376944 524418 376996 524424
rect 376942 523152 376998 523161
rect 376942 523087 376998 523096
rect 376956 523054 376984 523087
rect 376944 523048 376996 523054
rect 376944 522990 376996 522996
rect 376942 517984 376998 517993
rect 376942 517919 376998 517928
rect 376956 517546 376984 517919
rect 376944 517540 376996 517546
rect 376944 517482 376996 517488
rect 376942 515400 376998 515409
rect 376942 515335 376998 515344
rect 376956 514826 376984 515335
rect 376944 514820 376996 514826
rect 376944 514762 376996 514768
rect 376942 512816 376998 512825
rect 376942 512751 376998 512760
rect 376956 512038 376984 512751
rect 376944 512032 376996 512038
rect 376944 511974 376996 511980
rect 376942 510232 376998 510241
rect 376942 510167 376998 510176
rect 376956 509318 376984 510167
rect 376944 509312 376996 509318
rect 376944 509254 376996 509260
rect 268384 499520 268436 499526
rect 268384 499462 268436 499468
rect 267004 498160 267056 498166
rect 267004 498102 267056 498108
rect 377416 496806 377444 540903
rect 547156 538218 547184 552434
rect 551284 552424 551336 552430
rect 551284 552366 551336 552372
rect 548524 552356 548576 552362
rect 548524 552298 548576 552304
rect 547144 538212 547196 538218
rect 547144 538154 547196 538160
rect 377494 530768 377550 530777
rect 377494 530703 377550 530712
rect 377404 496800 377456 496806
rect 377404 496742 377456 496748
rect 264244 496732 264296 496738
rect 264244 496674 264296 496680
rect 377402 495000 377458 495009
rect 377402 494935 377458 494944
rect 377312 494760 377364 494766
rect 377312 494702 377364 494708
rect 262864 493944 262916 493950
rect 262864 493886 262916 493892
rect 376942 492416 376998 492425
rect 376942 492351 376998 492360
rect 260104 492040 260156 492046
rect 260104 491982 260156 491988
rect 376956 491366 376984 492351
rect 376944 491360 376996 491366
rect 376944 491302 376996 491308
rect 258724 491224 258776 491230
rect 258724 491166 258776 491172
rect 376942 489832 376998 489841
rect 376942 489767 376998 489776
rect 376956 488578 376984 489767
rect 376944 488572 376996 488578
rect 376944 488514 376996 488520
rect 255964 488504 256016 488510
rect 255964 488446 256016 488452
rect 376942 487248 376998 487257
rect 376942 487183 376944 487192
rect 376996 487183 376998 487192
rect 376944 487154 376996 487160
rect 253296 485648 253348 485654
rect 253296 485590 253348 485596
rect 377324 484362 377352 494702
rect 377312 484356 377364 484362
rect 377312 484298 377364 484304
rect 252468 482996 252520 483002
rect 252468 482938 252520 482944
rect 252376 482928 252428 482934
rect 252480 482905 252508 482938
rect 252376 482870 252428 482876
rect 252466 482896 252522 482905
rect 252388 482361 252416 482870
rect 252466 482831 252522 482840
rect 252374 482352 252430 482361
rect 252374 482287 252430 482296
rect 377218 482216 377274 482225
rect 377218 482151 377274 482160
rect 252468 480208 252520 480214
rect 252468 480150 252520 480156
rect 252480 480049 252508 480150
rect 252466 480040 252522 480049
rect 252466 479975 252522 479984
rect 377034 479632 377090 479641
rect 377034 479567 377090 479576
rect 252006 478544 252062 478553
rect 252006 478479 252062 478488
rect 251732 477430 251784 477436
rect 251914 477456 251970 477465
rect 251744 476785 251772 477430
rect 251914 477391 251970 477400
rect 376942 477048 376998 477057
rect 376942 476983 376998 476992
rect 251730 476776 251786 476785
rect 251730 476711 251786 476720
rect 376956 476134 376984 476983
rect 251916 476128 251968 476134
rect 251916 476070 251968 476076
rect 376944 476128 376996 476134
rect 376944 476070 376996 476076
rect 251928 473929 251956 476070
rect 252468 476060 252520 476066
rect 252468 476002 252520 476008
rect 252480 475697 252508 476002
rect 252466 475688 252522 475697
rect 252466 475623 252522 475632
rect 377048 474706 377076 479567
rect 377232 476066 377260 482151
rect 377416 480214 377444 494935
rect 377508 494018 377536 530703
rect 377586 520568 377642 520577
rect 377586 520503 377642 520512
rect 377496 494012 377548 494018
rect 377496 493954 377548 493960
rect 377600 489870 377628 520503
rect 377678 507784 377734 507793
rect 377678 507719 377734 507728
rect 377588 489864 377640 489870
rect 377588 489806 377640 489812
rect 377692 485790 377720 507719
rect 377770 505200 377826 505209
rect 377770 505135 377826 505144
rect 377784 494766 377812 505135
rect 377862 502616 377918 502625
rect 377862 502551 377918 502560
rect 377772 494760 377824 494766
rect 377772 494702 377824 494708
rect 377680 485784 377732 485790
rect 377680 485726 377732 485732
rect 377494 484664 377550 484673
rect 377494 484599 377550 484608
rect 377404 480208 377456 480214
rect 377404 480150 377456 480156
rect 377508 477494 377536 484599
rect 377876 483002 377904 502551
rect 377954 500032 378010 500041
rect 377954 499967 378010 499976
rect 377864 482996 377916 483002
rect 377864 482938 377916 482944
rect 377968 482934 377996 499967
rect 378046 497448 378102 497457
rect 378046 497383 378102 497392
rect 377956 482928 378008 482934
rect 377956 482870 378008 482876
rect 378060 481642 378088 497383
rect 378048 481636 378100 481642
rect 378048 481578 378100 481584
rect 377496 477488 377548 477494
rect 377496 477430 377548 477436
rect 377220 476060 377272 476066
rect 377220 476002 377272 476008
rect 252468 474700 252520 474706
rect 252468 474642 252520 474648
rect 377036 474700 377088 474706
rect 377036 474642 377088 474648
rect 252480 474473 252508 474642
rect 252466 474464 252522 474473
rect 252466 474399 252522 474408
rect 376942 474464 376998 474473
rect 376942 474399 376998 474408
rect 251914 473920 251970 473929
rect 251914 473855 251970 473864
rect 376956 473414 376984 474399
rect 251548 473408 251600 473414
rect 251548 473350 251600 473356
rect 376944 473408 376996 473414
rect 376944 473350 376996 473356
rect 251560 472977 251588 473350
rect 251546 472968 251602 472977
rect 251546 472903 251602 472912
rect 376942 471880 376998 471889
rect 376942 471815 376998 471824
rect 252466 471472 252522 471481
rect 252466 471407 252522 471416
rect 252480 471306 252508 471407
rect 376956 471306 376984 471815
rect 252468 471300 252520 471306
rect 252468 471242 252520 471248
rect 376944 471300 376996 471306
rect 376944 471242 376996 471248
rect 252466 470792 252522 470801
rect 252466 470727 252522 470736
rect 252480 470558 252508 470727
rect 252468 470552 252520 470558
rect 252468 470494 252520 470500
rect 376944 470552 376996 470558
rect 376944 470494 376996 470500
rect 376956 469305 376984 470494
rect 252466 469296 252522 469305
rect 252466 469231 252522 469240
rect 376942 469296 376998 469305
rect 376942 469231 376998 469240
rect 252374 468208 252430 468217
rect 252374 468143 252430 468152
rect 251546 467256 251602 467265
rect 251546 467191 251602 467200
rect 251270 464536 251326 464545
rect 251270 464471 251326 464480
rect 251284 463826 251312 464471
rect 251272 463820 251324 463826
rect 251272 463762 251324 463768
rect 251560 462330 251588 467191
rect 252282 465488 252338 465497
rect 252282 465423 252338 465432
rect 252190 463720 252246 463729
rect 252190 463655 252246 463664
rect 252006 462632 252062 462641
rect 252006 462567 252062 462576
rect 251548 462324 251600 462330
rect 251548 462266 251600 462272
rect 251914 461136 251970 461145
rect 251914 461071 251970 461080
rect 129752 460006 130686 460034
rect 131132 460006 132066 460034
rect 132512 460006 133538 460034
rect 133892 460006 134918 460034
rect 135272 460006 136390 460034
rect 136652 460006 137770 460034
rect 138032 460006 139242 460034
rect 139412 460006 140622 460034
rect 90364 457700 90416 457706
rect 90364 457642 90416 457648
rect 86224 457632 86276 457638
rect 86224 457574 86276 457580
rect 79324 457564 79376 457570
rect 79324 457506 79376 457512
rect 71320 392624 71372 392630
rect 71320 392566 71372 392572
rect 68744 391332 68796 391338
rect 68744 391274 68796 391280
rect 68756 386345 68784 391274
rect 71332 386345 71360 392566
rect 78496 386368 78548 386374
rect 68742 386336 68798 386345
rect 68742 386271 68798 386280
rect 71318 386336 71374 386345
rect 78494 386336 78496 386345
rect 78548 386336 78550 386345
rect 71318 386271 71374 386280
rect 73896 386300 73948 386306
rect 79336 386306 79364 457506
rect 80704 457496 80756 457502
rect 80704 457438 80756 457444
rect 80716 386374 80744 457438
rect 80704 386368 80756 386374
rect 80704 386310 80756 386316
rect 78494 386271 78550 386280
rect 79324 386300 79376 386306
rect 73896 386242 73948 386248
rect 79324 386242 79376 386248
rect 81072 386300 81124 386306
rect 81072 386242 81124 386248
rect 73908 385121 73936 386242
rect 77208 385892 77260 385898
rect 77208 385834 77260 385840
rect 77220 385121 77248 385834
rect 81084 385121 81112 386242
rect 86236 385150 86264 457574
rect 90376 386374 90404 457642
rect 126888 396908 126940 396914
rect 126888 396850 126940 396856
rect 124128 396840 124180 396846
rect 124128 396782 124180 396788
rect 121368 396772 121420 396778
rect 121368 396714 121420 396720
rect 118608 395684 118660 395690
rect 118608 395626 118660 395632
rect 117228 395616 117280 395622
rect 117228 395558 117280 395564
rect 114468 395548 114520 395554
rect 114468 395490 114520 395496
rect 111708 395480 111760 395486
rect 111708 395422 111760 395428
rect 108948 395412 109000 395418
rect 108948 395354 109000 395360
rect 106188 395344 106240 395350
rect 106188 395286 106240 395292
rect 104808 394256 104860 394262
rect 104808 394198 104860 394204
rect 102048 394188 102100 394194
rect 102048 394130 102100 394136
rect 99288 394120 99340 394126
rect 99288 394062 99340 394068
rect 96528 394052 96580 394058
rect 96528 393994 96580 394000
rect 93768 393984 93820 393990
rect 93768 393926 93820 393932
rect 89168 386368 89220 386374
rect 89166 386336 89168 386345
rect 90364 386368 90416 386374
rect 89220 386336 89222 386345
rect 93780 386345 93808 393926
rect 96540 386345 96568 393994
rect 99300 386345 99328 394062
rect 102060 386345 102088 394130
rect 90364 386310 90416 386316
rect 93766 386336 93822 386345
rect 89166 386271 89222 386280
rect 93766 386271 93822 386280
rect 96526 386336 96582 386345
rect 96526 386271 96582 386280
rect 99286 386336 99342 386345
rect 99286 386271 99342 386280
rect 102046 386336 102102 386345
rect 102046 386271 102102 386280
rect 86500 386232 86552 386238
rect 86500 386174 86552 386180
rect 83648 385144 83700 385150
rect 73894 385112 73950 385121
rect 73894 385047 73950 385056
rect 77206 385112 77262 385121
rect 77206 385047 77262 385056
rect 81070 385112 81126 385121
rect 81070 385047 81126 385056
rect 83646 385112 83648 385121
rect 86224 385144 86276 385150
rect 83700 385112 83702 385121
rect 86512 385121 86540 386174
rect 92112 386164 92164 386170
rect 92112 386106 92164 386112
rect 92124 385121 92152 386106
rect 104820 385257 104848 394198
rect 106200 386345 106228 395286
rect 108960 386345 108988 395354
rect 111720 386345 111748 395422
rect 106186 386336 106242 386345
rect 106186 386271 106242 386280
rect 108946 386336 109002 386345
rect 108946 386271 109002 386280
rect 111706 386336 111762 386345
rect 111706 386271 111762 386280
rect 104806 385248 104862 385257
rect 104806 385183 104862 385192
rect 114480 385121 114508 395490
rect 117240 386345 117268 395558
rect 118620 386345 118648 395626
rect 117226 386336 117282 386345
rect 117226 386271 117282 386280
rect 118606 386336 118662 386345
rect 118606 386271 118662 386280
rect 121380 385121 121408 396714
rect 124140 386345 124168 396782
rect 126900 386345 126928 396850
rect 129752 389842 129780 460006
rect 131132 389910 131160 460006
rect 132512 389978 132540 460006
rect 132500 389972 132552 389978
rect 132500 389914 132552 389920
rect 131120 389904 131172 389910
rect 131120 389846 131172 389852
rect 129740 389836 129792 389842
rect 129740 389778 129792 389784
rect 133696 386368 133748 386374
rect 124126 386336 124182 386345
rect 124126 386271 124182 386280
rect 126886 386336 126942 386345
rect 126886 386271 126942 386280
rect 133694 386336 133696 386345
rect 133748 386336 133750 386345
rect 133694 386271 133750 386280
rect 131028 386096 131080 386102
rect 131028 386038 131080 386044
rect 128636 385960 128688 385966
rect 128636 385902 128688 385908
rect 128648 385121 128676 385902
rect 131040 385121 131068 386038
rect 86224 385086 86276 385092
rect 86498 385112 86554 385121
rect 83646 385047 83702 385056
rect 86498 385047 86554 385056
rect 92110 385112 92166 385121
rect 92110 385047 92166 385056
rect 114466 385112 114522 385121
rect 114466 385047 114522 385056
rect 121366 385112 121422 385121
rect 121366 385047 121422 385056
rect 128634 385112 128690 385121
rect 128634 385047 128690 385056
rect 131026 385112 131082 385121
rect 131026 385047 131082 385056
rect 133892 384334 133920 460006
rect 134524 457768 134576 457774
rect 134524 457710 134576 457716
rect 134536 386374 134564 457710
rect 134524 386368 134576 386374
rect 134524 386310 134576 386316
rect 135272 384402 135300 460006
rect 136088 386028 136140 386034
rect 136088 385970 136140 385976
rect 136100 385121 136128 385970
rect 136086 385112 136142 385121
rect 136086 385047 136142 385056
rect 136652 384470 136680 460006
rect 138032 384538 138060 460006
rect 138480 386368 138532 386374
rect 138478 386336 138480 386345
rect 138532 386336 138534 386345
rect 138478 386271 138534 386280
rect 139412 384606 139440 460006
rect 142080 458046 142108 460020
rect 143460 458114 143488 460020
rect 143448 458108 143500 458114
rect 143448 458050 143500 458056
rect 142068 458040 142120 458046
rect 142068 457982 142120 457988
rect 140044 457836 140096 457842
rect 140044 457778 140096 457784
rect 140056 386374 140084 457778
rect 143448 397044 143500 397050
rect 143448 396986 143500 396992
rect 142068 396976 142120 396982
rect 142068 396918 142120 396924
rect 140044 386368 140096 386374
rect 142080 386345 142108 396918
rect 143460 386345 143488 396986
rect 144932 390114 144960 460020
rect 144920 390108 144972 390114
rect 144920 390050 144972 390056
rect 146312 387734 146340 460020
rect 147692 460006 147798 460034
rect 149072 460006 149178 460034
rect 150452 460006 150650 460034
rect 151832 460006 152030 460034
rect 153212 460006 153502 460034
rect 154592 460006 154882 460034
rect 155972 460006 156354 460034
rect 157352 460006 157734 460034
rect 158732 460006 159206 460034
rect 160112 460006 160678 460034
rect 161492 460006 162058 460034
rect 162872 460006 163530 460034
rect 164252 460006 164910 460034
rect 165632 460006 166382 460034
rect 167012 460006 167762 460034
rect 168392 460006 169234 460034
rect 169772 460006 170614 460034
rect 171152 460006 172086 460034
rect 172532 460006 173466 460034
rect 173912 460006 174938 460034
rect 175292 460006 176318 460034
rect 176672 460006 177790 460034
rect 178052 460006 179170 460034
rect 179432 460006 180642 460034
rect 180812 460006 182022 460034
rect 182192 460006 183494 460034
rect 183572 460006 184874 460034
rect 147692 391678 147720 460006
rect 149072 393038 149100 460006
rect 149060 393032 149112 393038
rect 149060 392974 149112 392980
rect 150452 392970 150480 460006
rect 150440 392964 150492 392970
rect 150440 392906 150492 392912
rect 151832 392902 151860 460006
rect 152464 457972 152516 457978
rect 152464 457914 152516 457920
rect 151820 392896 151872 392902
rect 151820 392838 151872 392844
rect 147680 391672 147732 391678
rect 147680 391614 147732 391620
rect 146300 387728 146352 387734
rect 146300 387670 146352 387676
rect 146208 386368 146260 386374
rect 140044 386310 140096 386316
rect 142066 386336 142122 386345
rect 142066 386271 142122 386280
rect 143446 386336 143502 386345
rect 146208 386310 146260 386316
rect 143446 386271 143502 386280
rect 146220 385121 146248 386310
rect 152476 385966 152504 457914
rect 153212 392834 153240 460006
rect 153200 392828 153252 392834
rect 153200 392770 153252 392776
rect 154592 392766 154620 460006
rect 155224 457904 155276 457910
rect 155224 457846 155276 457852
rect 154580 392760 154632 392766
rect 154580 392702 154632 392708
rect 155236 386374 155264 457846
rect 155972 392698 156000 460006
rect 157352 394330 157380 460006
rect 157340 394324 157392 394330
rect 157340 394266 157392 394272
rect 155960 392692 156012 392698
rect 155960 392634 156012 392640
rect 158732 391610 158760 460006
rect 158720 391604 158772 391610
rect 158720 391546 158772 391552
rect 160112 391474 160140 460006
rect 161492 391542 161520 460006
rect 161480 391536 161532 391542
rect 161480 391478 161532 391484
rect 160100 391468 160152 391474
rect 160100 391410 160152 391416
rect 162872 391406 162900 460006
rect 162860 391400 162912 391406
rect 162860 391342 162912 391348
rect 159824 390244 159876 390250
rect 159824 390186 159876 390192
rect 158536 390176 158588 390182
rect 158536 390118 158588 390124
rect 155224 386368 155276 386374
rect 158548 386345 158576 390118
rect 159836 386345 159864 390186
rect 164252 387666 164280 460006
rect 164240 387660 164292 387666
rect 164240 387602 164292 387608
rect 165632 387598 165660 460006
rect 165620 387592 165672 387598
rect 165620 387534 165672 387540
rect 167012 387530 167040 460006
rect 167000 387524 167052 387530
rect 167000 387466 167052 387472
rect 168392 387462 168420 460006
rect 168380 387456 168432 387462
rect 168380 387398 168432 387404
rect 169772 387394 169800 460006
rect 169760 387388 169812 387394
rect 169760 387330 169812 387336
rect 171152 387326 171180 460006
rect 171140 387320 171192 387326
rect 171140 387262 171192 387268
rect 172532 387258 172560 460006
rect 172520 387252 172572 387258
rect 172520 387194 172572 387200
rect 173912 387122 173940 460006
rect 175292 387190 175320 460006
rect 176672 388890 176700 460006
rect 176660 388884 176712 388890
rect 176660 388826 176712 388832
rect 178052 388822 178080 460006
rect 178040 388816 178092 388822
rect 178040 388758 178092 388764
rect 179432 388754 179460 460006
rect 179420 388748 179472 388754
rect 179420 388690 179472 388696
rect 180812 388686 180840 460006
rect 180800 388680 180852 388686
rect 180800 388622 180852 388628
rect 182192 388550 182220 460006
rect 183572 388618 183600 460006
rect 186332 390046 186360 460020
rect 186320 390040 186372 390046
rect 186320 389982 186372 389988
rect 183560 388612 183612 388618
rect 183560 388554 183612 388560
rect 182180 388544 182232 388550
rect 182180 388486 182232 388492
rect 187712 388482 187740 460020
rect 189092 460006 189198 460034
rect 190472 460006 190670 460034
rect 191852 460006 192050 460034
rect 193232 460006 193522 460034
rect 194612 460006 194902 460034
rect 195992 460006 196374 460034
rect 197372 460006 197754 460034
rect 198752 460006 199226 460034
rect 200132 460006 200606 460034
rect 201512 460006 202078 460034
rect 202892 460006 203458 460034
rect 204272 460006 204930 460034
rect 205652 460006 206310 460034
rect 189092 391270 189120 460006
rect 189080 391264 189132 391270
rect 189080 391206 189132 391212
rect 187700 388476 187752 388482
rect 187700 388418 187752 388424
rect 175280 387184 175332 387190
rect 175280 387126 175332 387132
rect 173900 387116 173952 387122
rect 173900 387058 173952 387064
rect 155224 386310 155276 386316
rect 158534 386336 158590 386345
rect 158534 386271 158590 386280
rect 159822 386336 159878 386345
rect 159822 386271 159878 386280
rect 152464 385960 152516 385966
rect 152464 385902 152516 385908
rect 146206 385112 146262 385121
rect 146206 385047 146262 385056
rect 170864 384668 170916 384674
rect 170864 384610 170916 384616
rect 177304 384668 177356 384674
rect 177304 384610 177356 384616
rect 139400 384600 139452 384606
rect 139400 384542 139452 384548
rect 138020 384532 138072 384538
rect 138020 384474 138072 384480
rect 136640 384464 136692 384470
rect 136640 384406 136692 384412
rect 135260 384396 135312 384402
rect 135260 384338 135312 384344
rect 133880 384328 133932 384334
rect 133880 384270 133932 384276
rect 170876 384169 170904 384610
rect 170862 384160 170918 384169
rect 170862 384095 170918 384104
rect 38290 336832 38346 336841
rect 38290 336767 38346 336776
rect 176660 336796 176712 336802
rect 38304 233918 38332 336767
rect 176660 336738 176712 336744
rect 38750 335608 38806 335617
rect 38750 335543 38806 335552
rect 38382 333160 38438 333169
rect 38382 333095 38438 333104
rect 38292 233912 38344 233918
rect 38292 233854 38344 233860
rect 38396 229809 38424 333095
rect 38566 332616 38622 332625
rect 38566 332551 38622 332560
rect 38474 309360 38530 309369
rect 38474 309295 38530 309304
rect 38382 229800 38438 229809
rect 38382 229735 38438 229744
rect 38488 161430 38516 309295
rect 38476 161424 38528 161430
rect 38476 161366 38528 161372
rect 38580 158846 38608 332551
rect 38658 327584 38714 327593
rect 38658 327519 38714 327528
rect 38672 158914 38700 327519
rect 38764 180810 38792 335543
rect 39026 330440 39082 330449
rect 39026 330375 39082 330384
rect 38842 329896 38898 329905
rect 38842 329831 38898 329840
rect 38856 234122 38884 329831
rect 38934 307864 38990 307873
rect 38934 307799 38990 307808
rect 38948 235618 38976 307799
rect 38936 235612 38988 235618
rect 38936 235554 38988 235560
rect 38844 234116 38896 234122
rect 38844 234058 38896 234064
rect 39040 234054 39068 330375
rect 39118 308408 39174 308417
rect 39118 308343 39174 308352
rect 39132 299470 39160 308343
rect 163226 299568 163282 299577
rect 163226 299503 163282 299512
rect 163410 299568 163466 299577
rect 163410 299503 163466 299512
rect 39120 299464 39172 299470
rect 39120 299406 39172 299412
rect 39948 299464 40000 299470
rect 39948 299406 40000 299412
rect 39028 234048 39080 234054
rect 39028 233990 39080 233996
rect 38752 180804 38804 180810
rect 38752 180746 38804 180752
rect 38660 158908 38712 158914
rect 38660 158850 38712 158856
rect 38568 158840 38620 158846
rect 38568 158782 38620 158788
rect 39960 158778 39988 299406
rect 163240 298926 163268 299503
rect 163228 298920 163280 298926
rect 163228 298862 163280 298868
rect 163424 298790 163452 299503
rect 163412 298784 163464 298790
rect 163412 298726 163464 298732
rect 56506 298072 56562 298081
rect 56506 298007 56562 298016
rect 57886 298072 57942 298081
rect 57886 298007 57942 298016
rect 59266 298072 59322 298081
rect 59266 298007 59322 298016
rect 60646 298072 60702 298081
rect 60646 298007 60702 298016
rect 62026 298072 62082 298081
rect 62026 298007 62082 298016
rect 63406 298072 63462 298081
rect 63406 298007 63462 298016
rect 64786 298072 64842 298081
rect 64786 298007 64842 298016
rect 66166 298072 66222 298081
rect 66166 298007 66222 298016
rect 67546 298072 67602 298081
rect 67546 298007 67602 298016
rect 68742 298072 68798 298081
rect 68742 298007 68798 298016
rect 70306 298072 70362 298081
rect 70306 298007 70362 298016
rect 71686 298072 71742 298081
rect 71686 298007 71742 298016
rect 73066 298072 73122 298081
rect 73066 298007 73122 298016
rect 74446 298072 74502 298081
rect 74446 298007 74502 298016
rect 75826 298072 75882 298081
rect 75826 298007 75882 298016
rect 77022 298072 77078 298081
rect 77022 298007 77078 298016
rect 78494 298072 78550 298081
rect 78494 298007 78550 298016
rect 79966 298072 80022 298081
rect 79966 298007 80022 298016
rect 80702 298072 80758 298081
rect 80702 298007 80758 298016
rect 81254 298072 81310 298081
rect 81254 298007 81310 298016
rect 82726 298072 82782 298081
rect 82726 298007 82782 298016
rect 83370 298072 83426 298081
rect 83370 298007 83426 298016
rect 84014 298072 84070 298081
rect 84014 298007 84070 298016
rect 85486 298072 85542 298081
rect 85486 298007 85542 298016
rect 86222 298072 86278 298081
rect 86222 298007 86278 298016
rect 86774 298072 86830 298081
rect 86774 298007 86830 298016
rect 88154 298072 88210 298081
rect 88154 298007 88210 298016
rect 89626 298072 89682 298081
rect 89626 298007 89682 298016
rect 91006 298072 91062 298081
rect 91006 298007 91062 298016
rect 92386 298072 92442 298081
rect 92386 298007 92442 298016
rect 93766 298072 93822 298081
rect 93766 298007 93822 298016
rect 95146 298072 95202 298081
rect 95146 298007 95202 298016
rect 96434 298072 96490 298081
rect 96434 298007 96490 298016
rect 97906 298072 97962 298081
rect 97906 298007 97962 298016
rect 99194 298072 99250 298081
rect 99194 298007 99250 298016
rect 102046 298072 102102 298081
rect 102046 298007 102102 298016
rect 106186 298072 106242 298081
rect 106186 298007 106242 298016
rect 108486 298072 108542 298081
rect 108486 298007 108542 298016
rect 111706 298072 111762 298081
rect 111706 298007 111762 298016
rect 114466 298072 114522 298081
rect 114466 298007 114522 298016
rect 115938 298072 115994 298081
rect 115938 298007 115994 298016
rect 117410 298072 117466 298081
rect 117410 298007 117466 298016
rect 121366 298072 121422 298081
rect 121366 298007 121422 298016
rect 124126 298072 124182 298081
rect 124126 298007 124182 298016
rect 125874 298072 125930 298081
rect 125874 298007 125930 298016
rect 129646 298072 129702 298081
rect 129646 298007 129702 298016
rect 133786 298072 133842 298081
rect 133786 298007 133842 298016
rect 136086 298072 136142 298081
rect 136086 298007 136088 298016
rect 56520 233986 56548 298007
rect 57900 234190 57928 298007
rect 57888 234184 57940 234190
rect 57888 234126 57940 234132
rect 56508 233980 56560 233986
rect 56508 233922 56560 233928
rect 39948 158772 40000 158778
rect 39948 158714 40000 158720
rect 59280 158506 59308 298007
rect 60554 297936 60610 297945
rect 60554 297871 60610 297880
rect 60568 231198 60596 297871
rect 60556 231192 60608 231198
rect 60556 231134 60608 231140
rect 60660 158710 60688 298007
rect 62040 172514 62068 298007
rect 62028 172508 62080 172514
rect 62028 172450 62080 172456
rect 63420 164218 63448 298007
rect 64800 229945 64828 298007
rect 66180 230081 66208 298007
rect 66166 230072 66222 230081
rect 66166 230007 66222 230016
rect 64786 229936 64842 229945
rect 64786 229871 64842 229880
rect 63408 164212 63460 164218
rect 63408 164154 63460 164160
rect 60648 158704 60700 158710
rect 60648 158646 60700 158652
rect 59268 158500 59320 158506
rect 59268 158442 59320 158448
rect 67560 158438 67588 298007
rect 68756 232694 68784 298007
rect 68834 297936 68890 297945
rect 68834 297871 68836 297880
rect 68888 297871 68890 297880
rect 69664 297900 69716 297906
rect 68836 297842 68888 297848
rect 69664 297842 69716 297848
rect 68834 297800 68890 297809
rect 68834 297735 68890 297744
rect 68848 232830 68876 297735
rect 68836 232824 68888 232830
rect 68836 232766 68888 232772
rect 68744 232688 68796 232694
rect 68744 232630 68796 232636
rect 69676 158574 69704 297842
rect 70320 239465 70348 298007
rect 70306 239456 70362 239465
rect 71700 239426 71728 298007
rect 73080 240854 73108 298007
rect 74354 297936 74410 297945
rect 74354 297871 74410 297880
rect 73068 240848 73120 240854
rect 73068 240790 73120 240796
rect 70306 239391 70362 239400
rect 71688 239420 71740 239426
rect 71688 239362 71740 239368
rect 74368 230217 74396 297871
rect 74354 230208 74410 230217
rect 74354 230143 74410 230152
rect 74460 169726 74488 298007
rect 75840 189038 75868 298007
rect 77036 233102 77064 298007
rect 77114 297936 77170 297945
rect 77114 297871 77170 297880
rect 77128 236706 77156 297871
rect 77206 297800 77262 297809
rect 77206 297735 77262 297744
rect 77220 297362 77248 297735
rect 77208 297356 77260 297362
rect 77208 297298 77260 297304
rect 77116 236700 77168 236706
rect 77116 236642 77168 236648
rect 77024 233096 77076 233102
rect 77024 233038 77076 233044
rect 75828 189032 75880 189038
rect 75828 188974 75880 188980
rect 78508 178022 78536 298007
rect 78586 297936 78642 297945
rect 78586 297871 78642 297880
rect 78496 178016 78548 178022
rect 78496 177958 78548 177964
rect 74448 169720 74500 169726
rect 74448 169662 74500 169668
rect 78600 159254 78628 297871
rect 79980 235550 80008 298007
rect 80716 296818 80744 298007
rect 80704 296812 80756 296818
rect 80704 296754 80756 296760
rect 79968 235544 80020 235550
rect 79968 235486 80020 235492
rect 81268 232898 81296 298007
rect 82740 236842 82768 298007
rect 83384 296886 83412 298007
rect 83372 296880 83424 296886
rect 83372 296822 83424 296828
rect 82728 236836 82780 236842
rect 82728 236778 82780 236784
rect 84028 236774 84056 298007
rect 84016 236768 84068 236774
rect 84016 236710 84068 236716
rect 81256 232892 81308 232898
rect 81256 232834 81308 232840
rect 85500 159322 85528 298007
rect 86236 296954 86264 298007
rect 86224 296948 86276 296954
rect 86224 296890 86276 296896
rect 85488 159316 85540 159322
rect 85488 159258 85540 159264
rect 78588 159248 78640 159254
rect 78588 159190 78640 159196
rect 86788 159186 86816 298007
rect 88168 186318 88196 298007
rect 88246 297936 88302 297945
rect 88246 297871 88302 297880
rect 88156 186312 88208 186318
rect 88156 186254 88208 186260
rect 86776 159180 86828 159186
rect 86776 159122 86828 159128
rect 88260 158982 88288 297871
rect 89640 238134 89668 298007
rect 90914 297936 90970 297945
rect 90914 297871 90970 297880
rect 89628 238128 89680 238134
rect 89628 238070 89680 238076
rect 90928 238066 90956 297871
rect 90916 238060 90968 238066
rect 90916 238002 90968 238008
rect 91020 231334 91048 298007
rect 92294 297936 92350 297945
rect 92294 297871 92350 297880
rect 91008 231328 91060 231334
rect 91008 231270 91060 231276
rect 92308 159118 92336 297871
rect 92296 159112 92348 159118
rect 92296 159054 92348 159060
rect 88248 158976 88300 158982
rect 88248 158918 88300 158924
rect 92400 158642 92428 298007
rect 93674 297936 93730 297945
rect 93674 297871 93730 297880
rect 93688 218006 93716 297871
rect 93676 218000 93728 218006
rect 93676 217942 93728 217948
rect 92388 158636 92440 158642
rect 92388 158578 92440 158584
rect 69664 158568 69716 158574
rect 69664 158510 69716 158516
rect 67548 158432 67600 158438
rect 67548 158374 67600 158380
rect 93780 157826 93808 298007
rect 95160 159050 95188 298007
rect 96448 229770 96476 298007
rect 96526 297936 96582 297945
rect 96526 297871 96582 297880
rect 96436 229764 96488 229770
rect 96436 229706 96488 229712
rect 96540 160478 96568 297871
rect 97920 223582 97948 298007
rect 99102 297936 99158 297945
rect 99102 297871 99158 297880
rect 99116 229838 99144 297871
rect 99208 229974 99236 298007
rect 99286 297800 99342 297809
rect 99286 297735 99342 297744
rect 99196 229968 99248 229974
rect 99196 229910 99248 229916
rect 99104 229832 99156 229838
rect 99104 229774 99156 229780
rect 97908 223576 97960 223582
rect 97908 223518 97960 223524
rect 96528 160472 96580 160478
rect 96528 160414 96580 160420
rect 95148 159044 95200 159050
rect 95148 158986 95200 158992
rect 99300 157894 99328 297735
rect 102060 158166 102088 298007
rect 104806 296848 104862 296857
rect 104806 296783 104862 296792
rect 102048 158160 102100 158166
rect 102048 158102 102100 158108
rect 104820 158098 104848 296783
rect 104808 158092 104860 158098
rect 104808 158034 104860 158040
rect 106200 158030 106228 298007
rect 108500 238754 108528 298007
rect 108580 297220 108632 297226
rect 108580 297162 108632 297168
rect 108408 238726 108528 238754
rect 108212 231464 108264 231470
rect 108212 231406 108264 231412
rect 107660 223576 107712 223582
rect 107658 223544 107660 223553
rect 107712 223544 107714 223553
rect 107658 223479 107714 223488
rect 108224 219434 108252 231406
rect 108304 231396 108356 231402
rect 108304 231338 108356 231344
rect 108316 229094 108344 231338
rect 108408 229906 108436 238726
rect 108488 231260 108540 231266
rect 108488 231202 108540 231208
rect 108396 229900 108448 229906
rect 108396 229842 108448 229848
rect 108316 229066 108436 229094
rect 108132 219406 108252 219434
rect 107660 218000 107712 218006
rect 107660 217942 107712 217948
rect 107672 217841 107700 217942
rect 107658 217832 107714 217841
rect 107658 217767 107714 217776
rect 108132 190454 108160 219406
rect 108132 190426 108252 190454
rect 107660 189032 107712 189038
rect 107660 188974 107712 188980
rect 107672 188873 107700 188974
rect 107658 188864 107714 188873
rect 107658 188799 107714 188808
rect 107660 186312 107712 186318
rect 107660 186254 107712 186260
rect 107672 186153 107700 186254
rect 107658 186144 107714 186153
rect 107658 186079 107714 186088
rect 107660 180804 107712 180810
rect 107660 180746 107712 180752
rect 107672 180713 107700 180746
rect 107658 180704 107714 180713
rect 107658 180639 107714 180648
rect 107660 178016 107712 178022
rect 107658 177984 107660 177993
rect 107712 177984 107714 177993
rect 107658 177919 107714 177928
rect 107660 172508 107712 172514
rect 107660 172450 107712 172456
rect 107672 172417 107700 172450
rect 107658 172408 107714 172417
rect 107658 172343 107714 172352
rect 107660 169720 107712 169726
rect 107658 169688 107660 169697
rect 107712 169688 107714 169697
rect 107658 169623 107714 169632
rect 108224 166977 108252 190426
rect 108408 175273 108436 229066
rect 108500 226273 108528 231202
rect 108486 226264 108542 226273
rect 108486 226199 108542 226208
rect 108592 215257 108620 297162
rect 108948 297152 109000 297158
rect 108948 297094 109000 297100
rect 108856 297084 108908 297090
rect 108856 297026 108908 297032
rect 108672 297016 108724 297022
rect 108672 296958 108724 296964
rect 108578 215248 108634 215257
rect 108578 215183 108634 215192
rect 108684 212537 108712 296958
rect 108764 296744 108816 296750
rect 108764 296686 108816 296692
rect 108670 212528 108726 212537
rect 108670 212463 108726 212472
rect 108776 206961 108804 296686
rect 108762 206952 108818 206961
rect 108762 206887 108818 206896
rect 108868 196897 108896 297026
rect 108854 196888 108910 196897
rect 108854 196823 108910 196832
rect 108960 183433 108988 297094
rect 109224 240916 109276 240922
rect 109224 240858 109276 240864
rect 109040 235476 109092 235482
rect 109040 235418 109092 235424
rect 109052 191457 109080 235418
rect 109132 235408 109184 235414
rect 109132 235350 109184 235356
rect 109144 194177 109172 235350
rect 109236 199617 109264 240858
rect 109592 240780 109644 240786
rect 109592 240722 109644 240728
rect 109316 235340 109368 235346
rect 109316 235282 109368 235288
rect 109328 202337 109356 235282
rect 109408 235272 109460 235278
rect 109408 235214 109460 235220
rect 109420 209681 109448 235214
rect 109500 231532 109552 231538
rect 109500 231474 109552 231480
rect 109406 209672 109462 209681
rect 109406 209607 109462 209616
rect 109512 204921 109540 231474
rect 109604 220493 109632 240722
rect 111340 235612 111392 235618
rect 111340 235554 111392 235560
rect 110328 231124 110380 231130
rect 110328 231066 110380 231072
rect 110340 228993 110368 231066
rect 111352 229922 111380 235554
rect 111720 232626 111748 298007
rect 111708 232620 111760 232626
rect 111708 232562 111760 232568
rect 114480 232558 114508 298007
rect 115388 233028 115440 233034
rect 115388 232970 115440 232976
rect 114468 232552 114520 232558
rect 114468 232494 114520 232500
rect 115400 229922 115428 232970
rect 115952 231538 115980 298007
rect 117424 296750 117452 298007
rect 117412 296744 117464 296750
rect 117412 296686 117464 296692
rect 118240 233980 118292 233986
rect 118240 233922 118292 233928
rect 115940 231532 115992 231538
rect 115940 231474 115992 231480
rect 111352 229894 111688 229922
rect 115092 229894 115428 229922
rect 118252 229922 118280 233922
rect 121380 231538 121408 298007
rect 121736 232688 121788 232694
rect 121736 232630 121788 232636
rect 121368 231532 121420 231538
rect 121368 231474 121420 231480
rect 121748 229922 121776 232630
rect 124140 231606 124168 298007
rect 125888 297226 125916 298007
rect 125876 297220 125928 297226
rect 125876 297162 125928 297168
rect 129660 296750 129688 298007
rect 129648 296744 129700 296750
rect 129648 296686 129700 296692
rect 132592 234184 132644 234190
rect 132592 234126 132644 234132
rect 129372 233980 129424 233986
rect 129372 233922 129424 233928
rect 125876 232960 125928 232966
rect 125876 232902 125928 232908
rect 124128 231600 124180 231606
rect 124128 231542 124180 231548
rect 125888 229922 125916 232902
rect 129384 229922 129412 233922
rect 118252 229894 118588 229922
rect 121748 229894 122084 229922
rect 125580 229894 125916 229922
rect 129076 229894 129412 229922
rect 132604 229786 132632 234126
rect 133800 231674 133828 298007
rect 136140 298007 136142 298016
rect 139306 298072 139362 298081
rect 141054 298072 141110 298081
rect 139306 298007 139362 298016
rect 140044 298036 140096 298042
rect 136088 297978 136140 297984
rect 137284 296744 137336 296750
rect 137284 296686 137336 296692
rect 136364 234184 136416 234190
rect 136364 234126 136416 234132
rect 133788 231668 133840 231674
rect 133788 231610 133840 231616
rect 136376 229922 136404 234126
rect 137296 232762 137324 296686
rect 137284 232756 137336 232762
rect 137284 232698 137336 232704
rect 139320 231742 139348 298007
rect 141054 298007 141110 298016
rect 146206 298072 146262 298081
rect 146206 298007 146262 298016
rect 140044 297978 140096 297984
rect 139400 234116 139452 234122
rect 139400 234058 139452 234064
rect 139308 231736 139360 231742
rect 139308 231678 139360 231684
rect 136068 229894 136404 229922
rect 139412 229922 139440 234058
rect 140056 232694 140084 297978
rect 141068 297226 141096 298007
rect 141056 297220 141108 297226
rect 141056 297162 141108 297168
rect 142712 233096 142764 233102
rect 142712 233038 142764 233044
rect 140044 232688 140096 232694
rect 140044 232630 140096 232636
rect 142724 229922 142752 233038
rect 146220 230450 146248 298007
rect 162124 297220 162176 297226
rect 162124 297162 162176 297168
rect 160100 242208 160152 242214
rect 160100 242150 160152 242156
rect 157248 236904 157300 236910
rect 157248 236846 157300 236852
rect 146300 234048 146352 234054
rect 146300 233990 146352 233996
rect 150256 234048 150308 234054
rect 150256 233990 150308 233996
rect 146208 230444 146260 230450
rect 146208 230386 146260 230392
rect 146312 229922 146340 233990
rect 150268 229922 150296 233990
rect 153200 232824 153252 232830
rect 153200 232766 153252 232772
rect 139412 229894 139564 229922
rect 142724 229894 143060 229922
rect 146312 229894 146556 229922
rect 149960 229894 150296 229922
rect 153212 229922 153240 232766
rect 157260 229922 157288 236846
rect 153212 229894 153456 229922
rect 156952 229894 157288 229922
rect 160112 229922 160140 242150
rect 162136 232830 162164 297162
rect 176672 248414 176700 336738
rect 177316 309126 177344 384610
rect 190472 379506 190500 460006
rect 191852 390250 191880 460006
rect 191840 390244 191892 390250
rect 191840 390186 191892 390192
rect 193232 390182 193260 460006
rect 193220 390176 193272 390182
rect 193220 390118 193272 390124
rect 178684 379500 178736 379506
rect 178684 379442 178736 379448
rect 190460 379500 190512 379506
rect 190460 379442 190512 379448
rect 178696 379273 178724 379442
rect 178682 379264 178738 379273
rect 178682 379199 178738 379208
rect 194612 320142 194640 460006
rect 178684 320136 178736 320142
rect 178684 320078 178736 320084
rect 194600 320136 194652 320142
rect 194600 320078 194652 320084
rect 178696 319433 178724 320078
rect 178682 319424 178738 319433
rect 178682 319359 178738 319368
rect 195992 318782 196020 460006
rect 178960 318776 179012 318782
rect 178960 318718 179012 318724
rect 195980 318776 196032 318782
rect 195980 318718 196032 318724
rect 178972 317801 179000 318718
rect 178958 317792 179014 317801
rect 178958 317727 179014 317736
rect 197372 317422 197400 460006
rect 178960 317416 179012 317422
rect 178960 317358 179012 317364
rect 197360 317416 197412 317422
rect 197360 317358 197412 317364
rect 178972 316441 179000 317358
rect 178958 316432 179014 316441
rect 178958 316367 179014 316376
rect 198752 315994 198780 460006
rect 178592 315988 178644 315994
rect 178592 315930 178644 315936
rect 198740 315988 198792 315994
rect 198740 315930 198792 315936
rect 178604 314945 178632 315930
rect 178590 314936 178646 314945
rect 178590 314871 178646 314880
rect 200132 314634 200160 460006
rect 178684 314628 178736 314634
rect 178684 314570 178736 314576
rect 200120 314628 200172 314634
rect 200120 314570 200172 314576
rect 178696 313721 178724 314570
rect 178682 313712 178738 313721
rect 178682 313647 178738 313656
rect 182824 309188 182876 309194
rect 182824 309130 182876 309136
rect 177304 309120 177356 309126
rect 177304 309062 177356 309068
rect 177316 299470 177344 309062
rect 177304 299464 177356 299470
rect 177304 299406 177356 299412
rect 176672 248386 177528 248414
rect 174728 237040 174780 237046
rect 174728 236982 174780 236988
rect 167736 236972 167788 236978
rect 167736 236914 167788 236920
rect 163596 232892 163648 232898
rect 163596 232834 163648 232840
rect 162124 232824 162176 232830
rect 162124 232766 162176 232772
rect 163608 229922 163636 232834
rect 167748 229922 167776 236914
rect 170956 234116 171008 234122
rect 170956 234058 171008 234064
rect 170968 229922 170996 234058
rect 174740 229922 174768 236982
rect 160112 229894 160448 229922
rect 163608 229894 163944 229922
rect 167440 229894 167776 229922
rect 170936 229894 170996 229922
rect 174432 229894 174768 229922
rect 177500 229922 177528 248386
rect 181076 233912 181128 233918
rect 181076 233854 181128 233860
rect 181088 229922 181116 233854
rect 182836 233034 182864 309130
rect 201512 298926 201540 460006
rect 201500 298920 201552 298926
rect 201500 298862 201552 298868
rect 202892 298790 202920 460006
rect 204272 391338 204300 460006
rect 205652 392630 205680 460006
rect 207768 457570 207796 460020
rect 208412 460006 209162 460034
rect 207756 457564 207808 457570
rect 207756 457506 207808 457512
rect 205640 392624 205692 392630
rect 205640 392566 205692 392572
rect 204260 391332 204312 391338
rect 204260 391274 204312 391280
rect 208412 385898 208440 460006
rect 210620 457502 210648 460020
rect 211172 460006 212014 460034
rect 210608 457496 210660 457502
rect 210608 457438 210660 457444
rect 211172 386306 211200 460006
rect 213472 457638 213500 460020
rect 213932 460006 214866 460034
rect 213460 457632 213512 457638
rect 213460 457574 213512 457580
rect 211160 386300 211212 386306
rect 211160 386242 211212 386248
rect 213932 386238 213960 460006
rect 216324 457706 216352 460020
rect 216692 460006 217718 460034
rect 218072 460006 219190 460034
rect 219452 460006 220662 460034
rect 220832 460006 222042 460034
rect 222212 460006 223514 460034
rect 223592 460006 224894 460034
rect 216312 457700 216364 457706
rect 216312 457642 216364 457648
rect 213920 386232 213972 386238
rect 213920 386174 213972 386180
rect 216692 386170 216720 460006
rect 218072 393990 218100 460006
rect 218704 458108 218756 458114
rect 218704 458050 218756 458056
rect 218060 393984 218112 393990
rect 218060 393926 218112 393932
rect 216680 386164 216732 386170
rect 216680 386106 216732 386112
rect 208400 385892 208452 385898
rect 208400 385834 208452 385840
rect 217876 384668 217928 384674
rect 217876 384610 217928 384616
rect 216678 336832 216734 336841
rect 216678 336767 216680 336776
rect 216732 336767 216734 336776
rect 216680 336738 216732 336744
rect 217322 335880 217378 335889
rect 217322 335815 217378 335824
rect 216678 309904 216734 309913
rect 216678 309839 216734 309848
rect 216692 309194 216720 309839
rect 216680 309188 216732 309194
rect 216680 309130 216732 309136
rect 216772 309120 216824 309126
rect 216772 309062 216824 309068
rect 216784 308417 216812 309062
rect 216770 308408 216826 308417
rect 216770 308343 216826 308352
rect 202880 298784 202932 298790
rect 202880 298726 202932 298732
rect 203524 297288 203576 297294
rect 203524 297230 203576 297236
rect 202144 297220 202196 297226
rect 202144 297162 202196 297168
rect 198740 295996 198792 296002
rect 198740 295938 198792 295944
rect 198752 248414 198780 295938
rect 198752 248386 198872 248414
rect 191840 240984 191892 240990
rect 191840 240926 191892 240932
rect 188620 235612 188672 235618
rect 188620 235554 188672 235560
rect 182824 233028 182876 233034
rect 182824 232970 182876 232976
rect 185216 233028 185268 233034
rect 185216 232970 185268 232976
rect 185228 229922 185256 232970
rect 188632 229922 188660 235554
rect 191852 229922 191880 240926
rect 194968 235544 195020 235550
rect 194968 235486 195020 235492
rect 177500 229894 177928 229922
rect 181088 229894 181424 229922
rect 184920 229894 185256 229922
rect 188324 229894 188660 229922
rect 191820 229894 191880 229922
rect 194980 229922 195008 235486
rect 194980 229894 195316 229922
rect 198844 229786 198872 248386
rect 202156 233034 202184 297162
rect 202144 233028 202196 233034
rect 202144 232970 202196 232976
rect 203536 232966 203564 297230
rect 205640 296064 205692 296070
rect 205640 296006 205692 296012
rect 203524 232960 203576 232966
rect 203524 232902 203576 232908
rect 202604 232892 202656 232898
rect 202604 232834 202656 232840
rect 202616 229922 202644 232834
rect 202308 229894 202644 229922
rect 205652 229922 205680 296006
rect 208952 236836 209004 236842
rect 208952 236778 209004 236784
rect 208964 229922 208992 236778
rect 216588 235544 216640 235550
rect 216588 235486 216640 235492
rect 213092 232960 213144 232966
rect 213092 232902 213144 232908
rect 213104 229922 213132 232902
rect 216600 229922 216628 235486
rect 217336 234122 217364 335815
rect 217506 329896 217562 329905
rect 217506 329831 217562 329840
rect 217520 234190 217548 329831
rect 217888 308417 217916 384610
rect 217966 333704 218022 333713
rect 217966 333639 218022 333648
rect 217874 308408 217930 308417
rect 217874 308343 217930 308352
rect 217874 308000 217930 308009
rect 217874 307935 217930 307944
rect 217508 234184 217560 234190
rect 217508 234126 217560 234132
rect 217324 234116 217376 234122
rect 217324 234058 217376 234064
rect 217888 230110 217916 307935
rect 217980 231810 218008 333639
rect 218716 298110 218744 458050
rect 218796 458040 218848 458046
rect 218796 457982 218848 457988
rect 218704 298104 218756 298110
rect 218704 298046 218756 298052
rect 218808 298042 218836 457982
rect 218888 457564 218940 457570
rect 218888 457506 218940 457512
rect 218900 386102 218928 457506
rect 219452 394058 219480 460006
rect 220084 457496 220136 457502
rect 220084 457438 220136 457444
rect 219440 394052 219492 394058
rect 219440 393994 219492 394000
rect 218888 386096 218940 386102
rect 218888 386038 218940 386044
rect 220096 386034 220124 457438
rect 220832 394126 220860 460006
rect 222212 394194 222240 460006
rect 223592 394262 223620 460006
rect 226352 395350 226380 460020
rect 227732 395418 227760 460020
rect 229112 460006 229218 460034
rect 230492 460006 230598 460034
rect 231872 460006 232070 460034
rect 233252 460006 233450 460034
rect 234632 460006 234922 460034
rect 236012 460006 236302 460034
rect 237392 460006 237774 460034
rect 229112 395486 229140 460006
rect 230492 395554 230520 460006
rect 231872 395622 231900 460006
rect 233252 395690 233280 460006
rect 234632 396778 234660 460006
rect 236012 396846 236040 460006
rect 237392 396914 237420 460006
rect 239140 457978 239168 460020
rect 239128 457972 239180 457978
rect 239128 457914 239180 457920
rect 240612 457570 240640 460020
rect 241992 457774 242020 460020
rect 241980 457768 242032 457774
rect 241980 457710 242032 457716
rect 240600 457564 240652 457570
rect 240600 457506 240652 457512
rect 243464 457502 243492 460020
rect 244844 457842 244872 460020
rect 245672 460006 246330 460034
rect 247052 460006 247710 460034
rect 244832 457836 244884 457842
rect 244832 457778 244884 457784
rect 243452 457496 243504 457502
rect 243452 457438 243504 457444
rect 245672 396982 245700 460006
rect 247052 397050 247080 460006
rect 249168 457910 249196 460020
rect 251822 459912 251878 459921
rect 251822 459847 251878 459856
rect 249156 457904 249208 457910
rect 249156 457846 249208 457852
rect 251836 441590 251864 459847
rect 251928 444378 251956 461071
rect 252020 449886 252048 462567
rect 252098 461680 252154 461689
rect 252098 461615 252154 461624
rect 252008 449880 252060 449886
rect 252008 449822 252060 449828
rect 252112 447098 252140 461615
rect 252204 452606 252232 463655
rect 252296 456754 252324 465423
rect 252388 465050 252416 468143
rect 252480 467838 252508 469231
rect 252468 467832 252520 467838
rect 252468 467774 252520 467780
rect 376944 467832 376996 467838
rect 376944 467774 376996 467780
rect 376956 466857 376984 467774
rect 376942 466848 376998 466857
rect 376942 466783 376998 466792
rect 252466 466576 252522 466585
rect 252466 466511 252522 466520
rect 252376 465044 252428 465050
rect 252376 464986 252428 464992
rect 252480 459542 252508 466511
rect 376944 465044 376996 465050
rect 376944 464986 376996 464992
rect 376956 464273 376984 464986
rect 376942 464264 376998 464273
rect 376942 464199 376998 464208
rect 253204 463820 253256 463826
rect 253204 463762 253256 463768
rect 252468 459536 252520 459542
rect 252468 459478 252520 459484
rect 252284 456748 252336 456754
rect 252284 456690 252336 456696
rect 253216 455394 253244 463762
rect 376944 462324 376996 462330
rect 376944 462266 376996 462272
rect 376956 461689 376984 462266
rect 376942 461680 376998 461689
rect 376942 461615 376998 461624
rect 376944 459536 376996 459542
rect 376944 459478 376996 459484
rect 376956 459105 376984 459478
rect 376942 459096 376998 459105
rect 376942 459031 376998 459040
rect 376944 456748 376996 456754
rect 376944 456690 376996 456696
rect 376956 456521 376984 456690
rect 376942 456512 376998 456521
rect 376942 456447 376998 456456
rect 253204 455388 253256 455394
rect 253204 455330 253256 455336
rect 376944 455388 376996 455394
rect 376944 455330 376996 455336
rect 376956 454073 376984 455330
rect 376942 454064 376998 454073
rect 376942 453999 376998 454008
rect 252192 452600 252244 452606
rect 252192 452542 252244 452548
rect 376852 452600 376904 452606
rect 376852 452542 376904 452548
rect 376864 451489 376892 452542
rect 376850 451480 376906 451489
rect 376850 451415 376906 451424
rect 376944 449880 376996 449886
rect 376944 449822 376996 449828
rect 376956 448905 376984 449822
rect 376942 448896 376998 448905
rect 376942 448831 376998 448840
rect 252100 447092 252152 447098
rect 252100 447034 252152 447040
rect 376944 447092 376996 447098
rect 376944 447034 376996 447040
rect 376956 446321 376984 447034
rect 376942 446312 376998 446321
rect 376942 446247 376998 446256
rect 251916 444372 251968 444378
rect 251916 444314 251968 444320
rect 376852 444372 376904 444378
rect 376852 444314 376904 444320
rect 376864 443737 376892 444314
rect 376850 443728 376906 443737
rect 376850 443663 376906 443672
rect 251824 441584 251876 441590
rect 251824 441526 251876 441532
rect 376944 441584 376996 441590
rect 376944 441526 376996 441532
rect 376956 441289 376984 441526
rect 376942 441280 376998 441289
rect 376942 441215 376998 441224
rect 379532 440014 380696 440042
rect 380912 440014 382076 440042
rect 382292 440014 383548 440042
rect 383672 440014 385020 440042
rect 386432 440014 386492 440042
rect 387812 440014 387964 440042
rect 389192 440014 389436 440042
rect 390572 440014 390908 440042
rect 391952 440014 392380 440042
rect 393516 440014 393852 440042
rect 394712 440014 395324 440042
rect 396092 440014 396796 440042
rect 397932 440014 398268 440042
rect 398852 440014 399740 440042
rect 400232 440014 401212 440042
rect 402348 440014 402684 440042
rect 402992 440014 404156 440042
rect 405292 440014 405628 440042
rect 405752 440014 407100 440042
rect 408512 440014 408572 440042
rect 409892 440014 410044 440042
rect 411272 440014 411516 440042
rect 412652 440014 412988 440042
rect 414032 440014 414460 440042
rect 415596 440014 415932 440042
rect 416792 440014 417404 440042
rect 418172 440014 418876 440042
rect 420012 440014 420348 440042
rect 420932 440014 421820 440042
rect 422956 440014 423292 440042
rect 423692 440014 424764 440042
rect 425072 440014 426236 440042
rect 427372 440014 427708 440042
rect 427832 440014 429180 440042
rect 430592 440014 430652 440042
rect 431972 440014 432124 440042
rect 433352 440014 433596 440042
rect 434732 440014 435068 440042
rect 436112 440014 436540 440042
rect 437492 440014 438012 440042
rect 438872 440014 439484 440042
rect 440252 440014 440956 440042
rect 441632 440014 442428 440042
rect 443012 440014 443900 440042
rect 445036 440014 445372 440042
rect 445772 440014 446844 440042
rect 447152 440014 448316 440042
rect 448532 440014 449788 440042
rect 449912 440014 451260 440042
rect 452672 440014 452732 440042
rect 454052 440014 454204 440042
rect 455432 440014 455676 440042
rect 456812 440014 457056 440042
rect 458192 440014 458528 440042
rect 459572 440014 460000 440042
rect 460952 440014 461472 440042
rect 462608 440014 462944 440042
rect 463712 440014 464416 440042
rect 465092 440014 465888 440042
rect 466472 440014 467360 440042
rect 467852 440014 468832 440042
rect 469968 440014 470304 440042
rect 470612 440014 471776 440042
rect 471992 440014 473248 440042
rect 474384 440014 474720 440042
rect 476132 440014 476192 440042
rect 477512 440014 477664 440042
rect 478892 440014 479136 440042
rect 480364 440014 480608 440042
rect 481652 440014 482080 440042
rect 483032 440014 483552 440042
rect 484412 440014 485024 440042
rect 485792 440014 486496 440042
rect 487632 440014 487968 440042
rect 488552 440014 489440 440042
rect 489932 440014 490912 440042
rect 492048 440014 492384 440042
rect 492692 440014 493856 440042
rect 494992 440014 495328 440042
rect 496464 440014 496800 440042
rect 498212 440014 498272 440042
rect 499592 440014 499744 440042
rect 500972 440014 501216 440042
rect 502352 440014 502688 440042
rect 503824 440014 504160 440042
rect 505296 440014 505632 440042
rect 506492 440014 507104 440042
rect 508240 440014 508576 440042
rect 509712 440014 510048 440042
rect 510632 440014 511520 440042
rect 512656 440014 512992 440042
rect 514128 440014 514464 440042
rect 514772 440014 515936 440042
rect 517072 440014 517408 440042
rect 518544 440014 518880 440042
rect 520292 440014 520352 440042
rect 521672 440014 521824 440042
rect 523052 440014 523296 440042
rect 524432 440014 524768 440042
rect 525904 440014 526240 440042
rect 527376 440014 527712 440042
rect 528848 440014 529184 440042
rect 358084 438320 358136 438326
rect 358084 438262 358136 438268
rect 247040 397044 247092 397050
rect 247040 396986 247092 396992
rect 245660 396976 245712 396982
rect 245660 396918 245712 396924
rect 237380 396908 237432 396914
rect 237380 396850 237432 396856
rect 236000 396840 236052 396846
rect 236000 396782 236052 396788
rect 234620 396772 234672 396778
rect 234620 396714 234672 396720
rect 233240 395684 233292 395690
rect 233240 395626 233292 395632
rect 231860 395616 231912 395622
rect 231860 395558 231912 395564
rect 230480 395548 230532 395554
rect 230480 395490 230532 395496
rect 229100 395480 229152 395486
rect 229100 395422 229152 395428
rect 227720 395412 227772 395418
rect 227720 395354 227772 395360
rect 226340 395344 226392 395350
rect 226340 395286 226392 395292
rect 270500 394324 270552 394330
rect 270500 394266 270552 394272
rect 223580 394256 223632 394262
rect 223580 394198 223632 394204
rect 222200 394188 222252 394194
rect 222200 394130 222252 394136
rect 220820 394120 220872 394126
rect 220820 394062 220872 394068
rect 255320 393032 255372 393038
rect 255320 392974 255372 392980
rect 252560 391672 252612 391678
rect 252560 391614 252612 391620
rect 248512 390108 248564 390114
rect 248512 390050 248564 390056
rect 248524 386345 248552 390050
rect 249800 387728 249852 387734
rect 249800 387670 249852 387676
rect 248510 386336 248566 386345
rect 248510 386271 248566 386280
rect 249812 386073 249840 387670
rect 252572 386345 252600 391614
rect 255332 386345 255360 392974
rect 258264 392964 258316 392970
rect 258264 392906 258316 392912
rect 258276 386345 258304 392906
rect 260840 392896 260892 392902
rect 260840 392838 260892 392844
rect 260852 386345 260880 392838
rect 263600 392828 263652 392834
rect 263600 392770 263652 392776
rect 263612 386345 263640 392770
rect 264980 392760 265032 392766
rect 264980 392702 265032 392708
rect 264992 386345 265020 392702
rect 268108 392692 268160 392698
rect 268108 392634 268160 392640
rect 268120 386345 268148 392634
rect 270512 386345 270540 394266
rect 273260 391604 273312 391610
rect 273260 391546 273312 391552
rect 273272 386345 273300 391546
rect 277952 391536 278004 391542
rect 277952 391478 278004 391484
rect 276020 391468 276072 391474
rect 276020 391410 276072 391416
rect 252558 386336 252614 386345
rect 252558 386271 252614 386280
rect 255318 386336 255374 386345
rect 255318 386271 255374 386280
rect 258262 386336 258318 386345
rect 258262 386271 258318 386280
rect 260838 386336 260894 386345
rect 260838 386271 260894 386280
rect 263598 386336 263654 386345
rect 263598 386271 263654 386280
rect 264978 386336 265034 386345
rect 264978 386271 265034 386280
rect 268106 386336 268162 386345
rect 268106 386271 268162 386280
rect 270498 386336 270554 386345
rect 270498 386271 270554 386280
rect 273258 386336 273314 386345
rect 273258 386271 273314 386280
rect 249798 386064 249854 386073
rect 220084 386028 220136 386034
rect 249798 385999 249854 386008
rect 220084 385970 220136 385976
rect 276032 385121 276060 391410
rect 277964 386345 277992 391478
rect 280160 391400 280212 391406
rect 280160 391342 280212 391348
rect 280172 386345 280200 391342
rect 325884 391264 325936 391270
rect 325884 391206 325936 391212
rect 320180 390040 320232 390046
rect 320180 389982 320232 389988
rect 305000 388884 305052 388890
rect 305000 388826 305052 388832
rect 282920 387660 282972 387666
rect 282920 387602 282972 387608
rect 277950 386336 278006 386345
rect 277950 386271 278006 386280
rect 280158 386336 280214 386345
rect 280158 386271 280214 386280
rect 282932 385121 282960 387602
rect 285680 387592 285732 387598
rect 285680 387534 285732 387540
rect 285692 386209 285720 387534
rect 288440 387524 288492 387530
rect 288440 387466 288492 387472
rect 288452 386345 288480 387466
rect 289820 387456 289872 387462
rect 289820 387398 289872 387404
rect 288438 386336 288494 386345
rect 288438 386271 288494 386280
rect 289832 386209 289860 387398
rect 292580 387388 292632 387394
rect 292580 387330 292632 387336
rect 285678 386200 285734 386209
rect 285678 386135 285734 386144
rect 289818 386200 289874 386209
rect 289818 386135 289874 386144
rect 292592 385121 292620 387330
rect 295340 387320 295392 387326
rect 295340 387262 295392 387268
rect 295352 386345 295380 387262
rect 298100 387252 298152 387258
rect 298100 387194 298152 387200
rect 295338 386336 295394 386345
rect 295338 386271 295394 386280
rect 298112 385937 298140 387194
rect 302240 387184 302292 387190
rect 302240 387126 302292 387132
rect 300860 387116 300912 387122
rect 300860 387058 300912 387064
rect 298098 385928 298154 385937
rect 298098 385863 298154 385872
rect 300872 385121 300900 387058
rect 302252 385937 302280 387126
rect 305012 386345 305040 388826
rect 307760 388816 307812 388822
rect 307760 388758 307812 388764
rect 304998 386336 305054 386345
rect 304998 386271 305054 386280
rect 302238 385928 302294 385937
rect 302238 385863 302294 385872
rect 307772 385121 307800 388758
rect 310520 388748 310572 388754
rect 310520 388690 310572 388696
rect 310532 386345 310560 388690
rect 313280 388680 313332 388686
rect 313280 388622 313332 388628
rect 313292 386345 313320 388622
rect 317420 388612 317472 388618
rect 317420 388554 317472 388560
rect 316040 388544 316092 388550
rect 316040 388486 316092 388492
rect 310518 386336 310574 386345
rect 310518 386271 310574 386280
rect 313278 386336 313334 386345
rect 313278 386271 313334 386280
rect 316052 386073 316080 388486
rect 317432 386345 317460 388554
rect 320192 386345 320220 389982
rect 322940 388476 322992 388482
rect 322940 388418 322992 388424
rect 322952 386345 322980 388418
rect 317418 386336 317474 386345
rect 317418 386271 317474 386280
rect 320178 386336 320234 386345
rect 320178 386271 320234 386280
rect 322938 386336 322994 386345
rect 322938 386271 322994 386280
rect 316038 386064 316094 386073
rect 316038 385999 316094 386008
rect 325896 385121 325924 391206
rect 338120 389972 338172 389978
rect 338120 389914 338172 389920
rect 338132 386345 338160 389914
rect 339500 389904 339552 389910
rect 339500 389846 339552 389852
rect 339512 386345 339540 389846
rect 338118 386336 338174 386345
rect 338118 386271 338174 386280
rect 339498 386336 339554 386345
rect 339498 386271 339554 386280
rect 351000 385688 351052 385694
rect 351000 385630 351052 385636
rect 351012 385121 351040 385630
rect 276018 385112 276074 385121
rect 276018 385047 276074 385056
rect 282918 385112 282974 385121
rect 282918 385047 282974 385056
rect 292578 385112 292634 385121
rect 292578 385047 292634 385056
rect 300858 385112 300914 385121
rect 300858 385047 300914 385056
rect 307758 385112 307814 385121
rect 307758 385047 307814 385056
rect 325882 385112 325938 385121
rect 325882 385047 325938 385056
rect 350998 385112 351054 385121
rect 350998 385047 351054 385056
rect 351012 384674 351040 385047
rect 351000 384668 351052 384674
rect 351000 384610 351052 384616
rect 343364 298104 343416 298110
rect 235998 298072 236054 298081
rect 218796 298036 218848 298042
rect 235998 298007 236054 298016
rect 238114 298072 238170 298081
rect 238114 298007 238170 298016
rect 242806 298072 242862 298081
rect 242806 298007 242862 298016
rect 247038 298072 247094 298081
rect 247038 298007 247094 298016
rect 248418 298072 248474 298081
rect 248418 298007 248474 298016
rect 249798 298072 249854 298081
rect 249798 298007 249854 298016
rect 251086 298072 251142 298081
rect 251086 298007 251142 298016
rect 251362 298072 251418 298081
rect 251362 298007 251418 298016
rect 251546 298072 251602 298081
rect 251546 298007 251602 298016
rect 252558 298072 252614 298081
rect 252558 298007 252614 298016
rect 258170 298072 258226 298081
rect 258170 298007 258226 298016
rect 259458 298072 259514 298081
rect 259458 298007 259514 298016
rect 260194 298072 260250 298081
rect 260194 298007 260250 298016
rect 261114 298072 261170 298081
rect 261114 298007 261170 298016
rect 263690 298072 263746 298081
rect 263690 298007 263746 298016
rect 265070 298072 265126 298081
rect 265070 298007 265126 298016
rect 265346 298072 265402 298081
rect 265346 298007 265402 298016
rect 266358 298072 266414 298081
rect 266358 298007 266414 298016
rect 267830 298072 267886 298081
rect 267830 298007 267886 298016
rect 269762 298072 269818 298081
rect 269762 298007 269818 298016
rect 270498 298072 270554 298081
rect 270498 298007 270554 298016
rect 271878 298072 271934 298081
rect 271878 298007 271934 298016
rect 273258 298072 273314 298081
rect 273258 298007 273314 298016
rect 274638 298072 274694 298081
rect 274638 298007 274694 298016
rect 276018 298072 276074 298081
rect 276018 298007 276074 298016
rect 276754 298072 276810 298081
rect 276754 298007 276810 298016
rect 277490 298072 277546 298081
rect 277490 298007 277546 298016
rect 278778 298072 278834 298081
rect 278778 298007 278834 298016
rect 280158 298072 280214 298081
rect 280158 298007 280214 298016
rect 282918 298072 282974 298081
rect 282918 298007 282974 298016
rect 285954 298072 286010 298081
rect 285954 298007 286010 298016
rect 287610 298072 287666 298081
rect 287610 298007 287666 298016
rect 290002 298072 290058 298081
rect 290002 298007 290058 298016
rect 292578 298072 292634 298081
rect 292578 298007 292634 298016
rect 295338 298072 295394 298081
rect 295338 298007 295394 298016
rect 298466 298072 298522 298081
rect 298466 298007 298522 298016
rect 300858 298072 300914 298081
rect 300858 298007 300914 298016
rect 302330 298072 302386 298081
rect 302330 298007 302386 298016
rect 305090 298072 305146 298081
rect 305090 298007 305146 298016
rect 308586 298072 308642 298081
rect 308586 298007 308642 298016
rect 310978 298072 311034 298081
rect 310978 298007 311034 298016
rect 313278 298072 313334 298081
rect 313278 298007 313334 298016
rect 315762 298072 315818 298081
rect 315762 298007 315818 298016
rect 317418 298072 317474 298081
rect 317418 298007 317474 298016
rect 320914 298072 320970 298081
rect 320914 298007 320970 298016
rect 322938 298072 322994 298081
rect 322938 298007 322994 298016
rect 325698 298072 325754 298081
rect 325698 298007 325754 298016
rect 343178 298072 343234 298081
rect 343178 298007 343180 298016
rect 218796 297978 218848 297984
rect 229836 238128 229888 238134
rect 229836 238070 229888 238076
rect 222936 236768 222988 236774
rect 222936 236710 222988 236716
rect 219624 232620 219676 232626
rect 219624 232562 219676 232568
rect 217968 231804 218020 231810
rect 217968 231746 218020 231752
rect 217876 230104 217928 230110
rect 217876 230046 217928 230052
rect 205652 229894 205804 229922
rect 208964 229894 209300 229922
rect 212796 229894 213132 229922
rect 216292 229894 216628 229922
rect 219636 229922 219664 232562
rect 222948 229922 222976 236710
rect 226340 232552 226392 232558
rect 226340 232494 226392 232500
rect 226352 229922 226380 232494
rect 229848 229922 229876 238070
rect 233332 238060 233384 238066
rect 233332 238002 233384 238008
rect 233344 229922 233372 238002
rect 236012 233986 236040 298007
rect 237286 297936 237342 297945
rect 237286 297871 237342 297880
rect 236000 233980 236052 233986
rect 236000 233922 236052 233928
rect 236828 232756 236880 232762
rect 236828 232698 236880 232704
rect 236840 229922 236868 232698
rect 237300 231062 237328 297871
rect 238128 297294 238156 298007
rect 238116 297288 238168 297294
rect 238116 297230 238168 297236
rect 240046 296848 240102 296857
rect 240046 296783 240102 296792
rect 237288 231056 237340 231062
rect 237288 230998 237340 231004
rect 240060 230994 240088 296783
rect 240968 236768 241020 236774
rect 240968 236710 241020 236716
rect 240048 230988 240100 230994
rect 240048 230930 240100 230936
rect 240980 229922 241008 236710
rect 242820 232762 242848 298007
rect 244188 236836 244240 236842
rect 244188 236778 244240 236784
rect 242808 232756 242860 232762
rect 242808 232698 242860 232704
rect 244200 229922 244228 236778
rect 247052 234054 247080 298007
rect 248326 297936 248382 297945
rect 248326 297871 248382 297880
rect 247040 234048 247092 234054
rect 247040 233990 247092 233996
rect 247316 232688 247368 232694
rect 247316 232630 247368 232636
rect 219636 229894 219788 229922
rect 222948 229894 223284 229922
rect 226352 229894 226688 229922
rect 229848 229894 230184 229922
rect 233344 229894 233680 229922
rect 236840 229894 237176 229922
rect 240672 229894 241008 229922
rect 244168 229894 244228 229922
rect 247328 229922 247356 232630
rect 248340 230042 248368 297871
rect 248432 236910 248460 298007
rect 249812 236978 249840 298007
rect 249800 236972 249852 236978
rect 249800 236914 249852 236920
rect 248420 236904 248472 236910
rect 248420 236846 248472 236852
rect 251100 232694 251128 298007
rect 251376 237046 251404 298007
rect 251560 297158 251588 298007
rect 251548 297152 251600 297158
rect 251548 297094 251600 297100
rect 251364 237040 251416 237046
rect 251364 236982 251416 236988
rect 251088 232688 251140 232694
rect 251088 232630 251140 232636
rect 251456 232552 251508 232558
rect 251456 232494 251508 232500
rect 248328 230036 248380 230042
rect 248328 229978 248380 229984
rect 251468 229922 251496 232494
rect 252572 231470 252600 298007
rect 256606 296984 256662 296993
rect 256606 296919 256662 296928
rect 255318 296848 255374 296857
rect 255318 296783 255374 296792
rect 255332 235482 255360 296783
rect 255320 235476 255372 235482
rect 255320 235418 255372 235424
rect 254952 232620 255004 232626
rect 254952 232562 255004 232568
rect 252560 231464 252612 231470
rect 252560 231406 252612 231412
rect 254964 229922 254992 232562
rect 256620 231470 256648 296919
rect 256698 296848 256754 296857
rect 256698 296783 256754 296792
rect 258078 296848 258134 296857
rect 258078 296783 258134 296792
rect 256712 235414 256740 296783
rect 256700 235408 256752 235414
rect 256700 235350 256752 235356
rect 256608 231464 256660 231470
rect 256608 231406 256660 231412
rect 258092 231402 258120 296783
rect 258184 235618 258212 298007
rect 258354 297800 258410 297809
rect 258354 297735 258410 297744
rect 258368 296041 258396 297735
rect 259472 297090 259500 298007
rect 259552 297356 259604 297362
rect 259552 297298 259604 297304
rect 259460 297084 259512 297090
rect 259460 297026 259512 297032
rect 259460 296948 259512 296954
rect 259460 296890 259512 296896
rect 258354 296032 258410 296041
rect 258354 295967 258410 295976
rect 258172 235612 258224 235618
rect 258172 235554 258224 235560
rect 258172 232824 258224 232830
rect 258172 232766 258224 232772
rect 258080 231396 258132 231402
rect 258080 231338 258132 231344
rect 258184 229922 258212 232766
rect 259368 230444 259420 230450
rect 259368 230386 259420 230392
rect 247328 229894 247664 229922
rect 251160 229894 251496 229922
rect 254656 229894 254992 229922
rect 258152 229894 258212 229922
rect 132572 229758 132632 229786
rect 198812 229758 198872 229786
rect 259380 229537 259408 230386
rect 259366 229528 259422 229537
rect 259366 229463 259422 229472
rect 110326 228984 110382 228993
rect 110326 228919 110382 228928
rect 109590 220484 109646 220493
rect 109590 220419 109646 220428
rect 109498 204912 109554 204921
rect 109498 204847 109554 204856
rect 109314 202328 109370 202337
rect 109314 202263 109370 202272
rect 109222 199608 109278 199617
rect 109222 199543 109278 199552
rect 109130 194168 109186 194177
rect 109130 194103 109186 194112
rect 259472 191593 259500 296890
rect 259564 202745 259592 297298
rect 259736 296880 259788 296886
rect 259736 296822 259788 296828
rect 259644 296812 259696 296818
rect 259644 296754 259696 296760
rect 259656 205601 259684 296754
rect 259748 209137 259776 296822
rect 260208 296002 260236 298007
rect 260930 296848 260986 296857
rect 260930 296783 260986 296792
rect 260196 295996 260248 296002
rect 260196 295938 260248 295944
rect 260944 242214 260972 296783
rect 261128 296070 261156 298007
rect 263598 297936 263654 297945
rect 263598 297871 263654 297880
rect 262218 296848 262274 296857
rect 262218 296783 262274 296792
rect 261116 296064 261168 296070
rect 261116 296006 261168 296012
rect 260932 242208 260984 242214
rect 260932 242150 260984 242156
rect 260196 240848 260248 240854
rect 260196 240790 260248 240796
rect 260104 239420 260156 239426
rect 260104 239362 260156 239368
rect 260012 230036 260064 230042
rect 260012 229978 260064 229984
rect 259920 229968 259972 229974
rect 259920 229910 259972 229916
rect 259828 229832 259880 229838
rect 259828 229774 259880 229780
rect 259840 226273 259868 229774
rect 259932 228041 259960 229910
rect 259918 228032 259974 228041
rect 259918 227967 259974 227976
rect 259826 226264 259882 226273
rect 259826 226199 259882 226208
rect 259828 224256 259880 224262
rect 259828 224198 259880 224204
rect 259734 209128 259790 209137
rect 259734 209063 259790 209072
rect 259642 205592 259698 205601
rect 259642 205527 259698 205536
rect 259550 202736 259606 202745
rect 259550 202671 259606 202680
rect 259458 191584 259514 191593
rect 259458 191519 259514 191528
rect 109038 191448 109094 191457
rect 109038 191383 109094 191392
rect 108946 183424 109002 183433
rect 108946 183359 109002 183368
rect 108394 175264 108450 175273
rect 108394 175199 108450 175208
rect 108210 166968 108266 166977
rect 108210 166903 108266 166912
rect 107660 164212 107712 164218
rect 107660 164154 107712 164160
rect 107672 164121 107700 164154
rect 107658 164112 107714 164121
rect 107658 164047 107714 164056
rect 259840 162761 259868 224198
rect 260024 222306 260052 229978
rect 259932 222278 260052 222306
rect 259932 165345 259960 222278
rect 260012 222216 260064 222222
rect 260012 222158 260064 222164
rect 260024 172417 260052 222158
rect 260116 187717 260144 239362
rect 260208 192613 260236 240790
rect 260288 236700 260340 236706
rect 260288 236642 260340 236648
rect 260300 198869 260328 236642
rect 262232 235550 262260 296783
rect 262220 235544 262272 235550
rect 262220 235486 262272 235492
rect 261116 232756 261168 232762
rect 261116 232698 261168 232704
rect 260840 232688 260892 232694
rect 260840 232630 260892 232636
rect 260472 231056 260524 231062
rect 260472 230998 260524 231004
rect 260484 224262 260512 230998
rect 260564 230988 260616 230994
rect 260564 230930 260616 230936
rect 260472 224256 260524 224262
rect 260472 224198 260524 224204
rect 260576 222222 260604 230930
rect 260564 222216 260616 222222
rect 260564 222158 260616 222164
rect 260286 198860 260342 198869
rect 260286 198795 260342 198804
rect 260194 192604 260250 192613
rect 260194 192539 260250 192548
rect 260102 187708 260158 187717
rect 260102 187643 260158 187652
rect 260010 172408 260066 172417
rect 260010 172343 260066 172352
rect 260852 169289 260880 232630
rect 261024 231192 261076 231198
rect 261024 231134 261076 231140
rect 261036 229094 261064 231134
rect 260944 229066 261064 229094
rect 260944 173913 260972 229066
rect 261128 224330 261156 232698
rect 262680 231804 262732 231810
rect 262680 231746 262732 231752
rect 261300 231532 261352 231538
rect 261300 231474 261352 231480
rect 261208 231464 261260 231470
rect 261208 231406 261260 231412
rect 261116 224324 261168 224330
rect 261116 224266 261168 224272
rect 261220 224210 261248 231406
rect 261036 224182 261248 224210
rect 261036 178809 261064 224182
rect 261116 224120 261168 224126
rect 261116 224062 261168 224068
rect 261128 180305 261156 224062
rect 261312 219434 261340 231474
rect 262404 231328 262456 231334
rect 262404 231270 262456 231276
rect 262312 224256 262364 224262
rect 262312 224198 262364 224204
rect 261220 219406 261340 219434
rect 261220 212265 261248 219406
rect 261206 212256 261262 212265
rect 261206 212191 261262 212200
rect 262220 189984 262272 189990
rect 262218 189952 262220 189961
rect 262272 189952 262274 189961
rect 262218 189887 262274 189896
rect 262324 182073 262352 224198
rect 262416 195945 262444 231270
rect 262588 229900 262640 229906
rect 262588 229842 262640 229848
rect 262496 229764 262548 229770
rect 262496 229706 262548 229712
rect 262508 201113 262536 229706
rect 262600 206961 262628 229842
rect 262692 224262 262720 231746
rect 262956 231736 263008 231742
rect 262956 231678 263008 231684
rect 262864 231668 262916 231674
rect 262864 231610 262916 231616
rect 262772 231600 262824 231606
rect 262772 231542 262824 231548
rect 262680 224256 262732 224262
rect 262680 224198 262732 224204
rect 262784 223922 262812 231542
rect 262772 223916 262824 223922
rect 262772 223858 262824 223864
rect 262876 223802 262904 231610
rect 262692 223774 262904 223802
rect 262692 220289 262720 223774
rect 262772 223712 262824 223718
rect 262968 223666 262996 231678
rect 263048 230104 263100 230110
rect 263048 230046 263100 230052
rect 262772 223654 262824 223660
rect 262678 220280 262734 220289
rect 262678 220215 262734 220224
rect 262784 219434 262812 223654
rect 262876 223638 262996 223666
rect 262876 221785 262904 223638
rect 262956 223576 263008 223582
rect 262956 223518 263008 223524
rect 262968 223145 262996 223518
rect 262954 223136 263010 223145
rect 262954 223071 263010 223080
rect 262862 221776 262918 221785
rect 262862 221711 262918 221720
rect 262692 219406 262812 219434
rect 262692 215257 262720 219406
rect 262678 215248 262734 215257
rect 262678 215183 262734 215192
rect 262586 206952 262642 206961
rect 262586 206887 262642 206896
rect 262494 201104 262550 201113
rect 262494 201039 262550 201048
rect 262402 195936 262458 195945
rect 262402 195871 262458 195880
rect 262310 182064 262366 182073
rect 262310 181999 262366 182008
rect 261114 180296 261170 180305
rect 261114 180231 261170 180240
rect 261022 178800 261078 178809
rect 261022 178735 261078 178744
rect 260930 173904 260986 173913
rect 260930 173839 260986 173848
rect 260838 169280 260894 169289
rect 260838 169215 260894 169224
rect 259918 165336 259974 165345
rect 259918 165271 259974 165280
rect 259826 162752 259882 162761
rect 259826 162687 259882 162696
rect 107660 161424 107712 161430
rect 107658 161392 107660 161401
rect 107712 161392 107714 161401
rect 107658 161327 107714 161336
rect 263060 161129 263088 230046
rect 263508 224936 263560 224942
rect 263508 224878 263560 224884
rect 263520 224641 263548 224878
rect 263506 224632 263562 224641
rect 263506 224567 263562 224576
rect 263508 218000 263560 218006
rect 263506 217968 263508 217977
rect 263560 217968 263562 217977
rect 263506 217903 263562 217912
rect 263508 216640 263560 216646
rect 263508 216582 263560 216588
rect 263520 216481 263548 216582
rect 263506 216472 263562 216481
rect 263506 216407 263562 216416
rect 263508 213920 263560 213926
rect 263508 213862 263560 213868
rect 263520 213625 263548 213862
rect 263506 213616 263562 213625
rect 263506 213551 263562 213560
rect 263508 211132 263560 211138
rect 263508 211074 263560 211080
rect 263520 210633 263548 211074
rect 263506 210624 263562 210633
rect 263506 210559 263562 210568
rect 263508 204264 263560 204270
rect 263508 204206 263560 204212
rect 263520 203969 263548 204206
rect 263506 203960 263562 203969
rect 263506 203895 263562 203904
rect 263046 161120 263102 161129
rect 263046 161055 263102 161064
rect 110604 160472 110656 160478
rect 216770 160440 216826 160449
rect 110604 160414 110656 160420
rect 110492 160126 110552 160154
rect 110420 159384 110472 159390
rect 110420 159326 110472 159332
rect 110432 158778 110460 159326
rect 110420 158772 110472 158778
rect 110420 158714 110472 158720
rect 106188 158024 106240 158030
rect 106188 157966 106240 157972
rect 99288 157888 99340 157894
rect 99288 157830 99340 157836
rect 93768 157820 93820 157826
rect 93768 157762 93820 157768
rect 106280 38344 106332 38350
rect 106280 38286 106332 38292
rect 99380 38276 99432 38282
rect 99380 38218 99432 38224
rect 50344 38208 50396 38214
rect 50344 38150 50396 38156
rect 35164 38072 35216 38078
rect 35164 38014 35216 38020
rect 22744 38004 22796 38010
rect 22744 37946 22796 37952
rect 10324 37936 10376 37942
rect 10324 37878 10376 37884
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 572 9376 624 9382
rect 572 9318 624 9324
rect 584 480 612 9318
rect 1676 9240 1728 9246
rect 1676 9182 1728 9188
rect 1688 480 1716 9182
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 480 2912 8910
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 480 4108 6122
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 480 5304 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 8978
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8772 480 8800 6190
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 17206
rect 10336 3534 10364 37878
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13832 16574 13860 19926
rect 13832 16546 14320 16574
rect 13544 13116 13596 13122
rect 13544 13058 13596 13064
rect 11888 10328 11940 10334
rect 11888 10270 11940 10276
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 10270
rect 13556 480 13584 13058
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17052 480 17080 11698
rect 18236 7608 18288 7614
rect 18236 7550 18288 7556
rect 18248 480 18276 7550
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19444 480 19472 3130
rect 21836 480 21864 11766
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 15846
rect 22756 3194 22784 37946
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 27712 15972 27764 15978
rect 27712 15914 27764 15920
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 24228 480 24256 3470
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 13126
rect 27724 480 27752 15914
rect 30104 6520 30156 6526
rect 30104 6462 30156 6468
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30116 480 30144 6462
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 15982
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 32416 480 32444 3538
rect 33612 480 33640 13262
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 16050
rect 35176 3398 35204 38014
rect 45560 21412 45612 21418
rect 45560 21354 45612 21360
rect 44180 17604 44232 17610
rect 44180 17546 44232 17552
rect 41420 17536 41472 17542
rect 41420 17478 41472 17484
rect 41432 16574 41460 17478
rect 44192 16574 44220 17546
rect 45572 16574 45600 21354
rect 49700 17332 49752 17338
rect 49700 17274 49752 17280
rect 49712 16574 49740 17274
rect 41432 16546 41920 16574
rect 44192 16546 45048 16574
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 38384 16176 38436 16182
rect 38384 16118 38436 16124
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36004 480 36032 3674
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 13330
rect 38396 480 38424 16118
rect 40684 6588 40736 6594
rect 40684 6530 40736 6536
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39592 480 39620 3606
rect 40696 480 40724 6530
rect 41892 480 41920 16546
rect 44272 6656 44324 6662
rect 44272 6598 44324 6604
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 43088 480 43116 3742
rect 44284 480 44312 6598
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 47860 9104 47912 9110
rect 47860 9046 47912 9052
rect 47872 480 47900 9046
rect 48964 6316 49016 6322
rect 48964 6258 49016 6264
rect 48976 480 49004 6258
rect 50172 480 50200 16546
rect 50356 3738 50384 38150
rect 51724 38140 51776 38146
rect 51724 38082 51776 38088
rect 51356 9172 51408 9178
rect 51356 9114 51408 9120
rect 50344 3732 50396 3738
rect 50344 3674 50396 3680
rect 51368 480 51396 9114
rect 51736 3806 51764 38082
rect 95240 20324 95292 20330
rect 95240 20266 95292 20272
rect 92480 20256 92532 20262
rect 92480 20198 92532 20204
rect 88340 20188 88392 20194
rect 88340 20130 88392 20136
rect 85580 20120 85632 20126
rect 85580 20062 85632 20068
rect 81440 20052 81492 20058
rect 81440 19994 81492 20000
rect 77300 18964 77352 18970
rect 77300 18906 77352 18912
rect 74540 18896 74592 18902
rect 74540 18838 74592 18844
rect 70400 18828 70452 18834
rect 70400 18770 70452 18776
rect 67640 18760 67692 18766
rect 67640 18702 67692 18708
rect 63500 18692 63552 18698
rect 63500 18634 63552 18640
rect 60740 18624 60792 18630
rect 60740 18566 60792 18572
rect 56600 17468 56652 17474
rect 56600 17410 56652 17416
rect 52460 17400 52512 17406
rect 52460 17342 52512 17348
rect 52472 16574 52500 17342
rect 56612 16574 56640 17410
rect 60752 16574 60780 18566
rect 63512 16574 63540 18634
rect 52472 16546 53328 16574
rect 56612 16546 56824 16574
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 52552 6384 52604 6390
rect 52552 6326 52604 6332
rect 51724 3800 51776 3806
rect 51724 3742 51776 3748
rect 52564 480 52592 6326
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54944 10396 54996 10402
rect 54944 10338 54996 10344
rect 54956 480 54984 10338
rect 56048 6452 56100 6458
rect 56048 6394 56100 6400
rect 56060 480 56088 6394
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 59360 13252 59412 13258
rect 59360 13194 59412 13200
rect 58440 10464 58492 10470
rect 58440 10406 58492 10412
rect 58452 480 58480 10406
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13194
rect 60844 480 60872 16546
rect 63224 14476 63276 14482
rect 63224 14418 63276 14424
rect 61568 10532 61620 10538
rect 61568 10474 61620 10480
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 10474
rect 63236 480 63264 14418
rect 64340 480 64368 16546
rect 66720 14544 66772 14550
rect 66720 14486 66772 14492
rect 65064 10600 65116 10606
rect 65064 10542 65116 10548
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 10542
rect 66732 480 66760 14486
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 18702
rect 70412 16574 70440 18770
rect 74552 16574 74580 18838
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 69020 14612 69072 14618
rect 69020 14554 69072 14560
rect 69032 3398 69060 14554
rect 69112 10668 69164 10674
rect 69112 10610 69164 10616
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 69124 480 69152 10610
rect 69940 3392 69992 3398
rect 69940 3334 69992 3340
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3334
rect 71516 480 71544 16546
rect 73344 14680 73396 14686
rect 73344 14622 73396 14628
rect 72608 4820 72660 4826
rect 72608 4762 72660 4768
rect 72620 480 72648 4762
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 14622
rect 75012 480 75040 16546
rect 76196 4888 76248 4894
rect 76196 4830 76248 4836
rect 76208 480 76236 4830
rect 77312 3398 77340 18906
rect 81452 16574 81480 19994
rect 85592 16574 85620 20062
rect 88352 16574 88380 20130
rect 81452 16546 81664 16574
rect 85592 16546 85712 16574
rect 88352 16546 89208 16574
rect 80888 14816 80940 14822
rect 80888 14758 80940 14764
rect 77392 14748 77444 14754
rect 77392 14690 77444 14696
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 14690
rect 79692 4956 79744 4962
rect 79692 4898 79744 4904
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 79704 480 79732 4898
rect 80900 480 80928 14758
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 84200 16244 84252 16250
rect 84200 16186 84252 16192
rect 83280 5024 83332 5030
rect 83280 4966 83332 4972
rect 83292 480 83320 4966
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 16186
rect 85684 480 85712 16546
rect 87972 7676 88024 7682
rect 87972 7618 88024 7624
rect 86868 5092 86920 5098
rect 86868 5034 86920 5040
rect 86880 480 86908 5034
rect 87984 480 88012 7618
rect 89180 480 89208 16546
rect 91560 7744 91612 7750
rect 91560 7686 91612 7692
rect 90364 5160 90416 5166
rect 90364 5102 90416 5108
rect 90376 480 90404 5102
rect 91572 480 91600 7686
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 20198
rect 95252 16574 95280 20266
rect 99392 16574 99420 38218
rect 102140 21480 102192 21486
rect 102140 21422 102192 21428
rect 95252 16546 95832 16574
rect 99392 16546 99880 16574
rect 93952 11892 94004 11898
rect 93952 11834 94004 11840
rect 93964 480 93992 11834
rect 95148 7812 95200 7818
rect 95148 7754 95200 7760
rect 95160 480 95188 7754
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 97448 11960 97500 11966
rect 97448 11902 97500 11908
rect 97460 480 97488 11902
rect 98644 7880 98696 7886
rect 98644 7822 98696 7828
rect 98656 480 98684 7822
rect 99852 480 99880 16546
rect 101036 5228 101088 5234
rect 101036 5170 101088 5176
rect 101048 480 101076 5170
rect 102152 3398 102180 21422
rect 106292 16574 106320 38286
rect 106292 16546 106504 16574
rect 104072 12028 104124 12034
rect 104072 11970 104124 11976
rect 102232 7948 102284 7954
rect 102232 7890 102284 7896
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 7890
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 11970
rect 105728 8016 105780 8022
rect 105728 7958 105780 7964
rect 105740 480 105768 7958
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 110432 9382 110460 158714
rect 110524 118658 110552 160126
rect 110616 158370 110644 160414
rect 216568 160398 216770 160426
rect 218886 160440 218942 160449
rect 218592 160398 218886 160426
rect 216770 160375 216826 160384
rect 218886 160375 218942 160384
rect 161460 160262 161704 160290
rect 111168 160126 111504 160154
rect 111812 160126 112516 160154
rect 113192 160126 113528 160154
rect 114540 160126 114692 160154
rect 111168 159390 111196 160126
rect 111156 159384 111208 159390
rect 111156 159326 111208 159332
rect 110604 158364 110656 158370
rect 110604 158306 110656 158312
rect 111812 120086 111840 160126
rect 113192 158778 113220 160126
rect 113180 158772 113232 158778
rect 113180 158714 113232 158720
rect 111800 120080 111852 120086
rect 111800 120022 111852 120028
rect 110512 118652 110564 118658
rect 110512 118594 110564 118600
rect 110512 21548 110564 21554
rect 110512 21490 110564 21496
rect 110420 9376 110472 9382
rect 110420 9318 110472 9324
rect 108120 9308 108172 9314
rect 108120 9250 108172 9256
rect 108132 480 108160 9250
rect 109316 8084 109368 8090
rect 109316 8026 109368 8032
rect 109328 480 109356 8026
rect 110524 480 110552 21490
rect 111616 12096 111668 12102
rect 111616 12038 111668 12044
rect 111628 480 111656 12038
rect 113192 9246 113220 158714
rect 114560 155984 114612 155990
rect 114560 155926 114612 155932
rect 114572 117298 114600 155926
rect 114664 118590 114692 160126
rect 115216 160126 115552 160154
rect 115952 160126 116564 160154
rect 117424 160126 117576 160154
rect 118252 160126 118588 160154
rect 118712 160126 119600 160154
rect 120092 160126 120612 160154
rect 121624 160126 121684 160154
rect 115216 155990 115244 160126
rect 115204 155984 115256 155990
rect 115204 155926 115256 155932
rect 114652 118584 114704 118590
rect 114652 118526 114704 118532
rect 114560 117292 114612 117298
rect 114560 117234 114612 117240
rect 115952 41410 115980 160126
rect 117320 155984 117372 155990
rect 117320 155926 117372 155932
rect 117332 66230 117360 155926
rect 117424 92478 117452 160126
rect 118252 155990 118280 160126
rect 118240 155984 118292 155990
rect 118240 155926 118292 155932
rect 117412 92472 117464 92478
rect 117412 92414 117464 92420
rect 117320 66224 117372 66230
rect 117320 66166 117372 66172
rect 115940 41404 115992 41410
rect 115940 41346 115992 41352
rect 118712 41342 118740 160126
rect 120092 92410 120120 160126
rect 121460 155984 121512 155990
rect 121460 155926 121512 155932
rect 120080 92404 120132 92410
rect 120080 92346 120132 92352
rect 121472 42770 121500 155926
rect 121656 142154 121684 160126
rect 122392 160126 122728 160154
rect 122852 160126 123740 160154
rect 124232 160126 124752 160154
rect 125612 160126 125764 160154
rect 126256 160126 126776 160154
rect 126992 160126 127788 160154
rect 128372 160126 128800 160154
rect 129812 160126 129872 160154
rect 122392 155990 122420 160126
rect 122380 155984 122432 155990
rect 122380 155926 122432 155932
rect 121564 142126 121684 142154
rect 121564 67590 121592 142126
rect 122852 93838 122880 160126
rect 122840 93832 122892 93838
rect 122840 93774 122892 93780
rect 121552 67584 121604 67590
rect 121552 67526 121604 67532
rect 124232 67522 124260 160126
rect 124220 67516 124272 67522
rect 124220 67458 124272 67464
rect 121460 42764 121512 42770
rect 121460 42706 121512 42712
rect 125612 42702 125640 160126
rect 126256 142154 126284 160126
rect 125704 142126 126284 142154
rect 125704 93770 125732 142126
rect 125692 93764 125744 93770
rect 125692 93706 125744 93712
rect 126992 69018 127020 160126
rect 126980 69012 127032 69018
rect 126980 68954 127032 68960
rect 128372 44130 128400 160126
rect 129740 155984 129792 155990
rect 129740 155926 129792 155932
rect 129752 70378 129780 155926
rect 129844 95198 129872 160126
rect 130488 160126 130824 160154
rect 131132 160126 131836 160154
rect 132512 160126 132848 160154
rect 133952 160126 134012 160154
rect 130488 155990 130516 160126
rect 130476 155984 130528 155990
rect 130476 155926 130528 155932
rect 129832 95192 129884 95198
rect 129832 95134 129884 95140
rect 129740 70372 129792 70378
rect 129740 70314 129792 70320
rect 131132 45558 131160 160126
rect 132512 96626 132540 160126
rect 133880 155984 133932 155990
rect 133880 155926 133932 155932
rect 132500 96620 132552 96626
rect 132500 96562 132552 96568
rect 131120 45552 131172 45558
rect 131120 45494 131172 45500
rect 133892 45490 133920 155926
rect 133984 70310 134012 160126
rect 134628 160126 134964 160154
rect 135272 160126 135976 160154
rect 136652 160126 136988 160154
rect 138000 160126 138060 160154
rect 134628 155990 134656 160126
rect 134616 155984 134668 155990
rect 134616 155926 134668 155932
rect 135272 96558 135300 160126
rect 135260 96552 135312 96558
rect 135260 96494 135312 96500
rect 136652 71738 136680 160126
rect 136640 71732 136692 71738
rect 136640 71674 136692 71680
rect 133972 70304 134024 70310
rect 133972 70246 134024 70252
rect 138032 46918 138060 160126
rect 138124 160126 139012 160154
rect 139412 160126 140024 160154
rect 140792 160126 141036 160154
rect 141160 160126 142048 160154
rect 142172 160126 143060 160154
rect 143552 160126 144072 160154
rect 145024 160126 145176 160154
rect 145852 160126 146188 160154
rect 146312 160126 147200 160154
rect 147692 160126 148212 160154
rect 149224 160126 149284 160154
rect 138124 97986 138152 160126
rect 138112 97980 138164 97986
rect 138112 97922 138164 97928
rect 139412 71670 139440 160126
rect 139400 71664 139452 71670
rect 139400 71606 139452 71612
rect 138020 46912 138072 46918
rect 138020 46854 138072 46860
rect 140792 46850 140820 160126
rect 141160 142154 141188 160126
rect 140884 142126 141188 142154
rect 140884 97918 140912 142126
rect 140872 97912 140924 97918
rect 140872 97854 140924 97860
rect 142172 73166 142200 160126
rect 142160 73160 142212 73166
rect 142160 73102 142212 73108
rect 143552 48278 143580 160126
rect 144920 155984 144972 155990
rect 144920 155926 144972 155932
rect 144932 73098 144960 155926
rect 145024 99346 145052 160126
rect 145852 155990 145880 160126
rect 145840 155984 145892 155990
rect 145840 155926 145892 155932
rect 145012 99340 145064 99346
rect 145012 99282 145064 99288
rect 144920 73092 144972 73098
rect 144920 73034 144972 73040
rect 143540 48272 143592 48278
rect 143540 48214 143592 48220
rect 146312 48210 146340 160126
rect 147692 100706 147720 160126
rect 149060 155984 149112 155990
rect 149060 155926 149112 155932
rect 147680 100700 147732 100706
rect 147680 100642 147732 100648
rect 149072 49706 149100 155926
rect 149256 142154 149284 160126
rect 149900 160126 150236 160154
rect 150452 160126 151248 160154
rect 151832 160126 152260 160154
rect 153272 160126 153332 160154
rect 149900 155990 149928 160126
rect 149888 155984 149940 155990
rect 149888 155926 149940 155932
rect 149164 142126 149284 142154
rect 149164 74526 149192 142126
rect 150452 100638 150480 160126
rect 150440 100632 150492 100638
rect 150440 100574 150492 100580
rect 151832 75886 151860 160126
rect 153304 155938 153332 160126
rect 153212 155910 153332 155938
rect 153396 160126 154284 160154
rect 154592 160126 155296 160154
rect 155972 160126 156308 160154
rect 157412 160126 157472 160154
rect 151820 75880 151872 75886
rect 151820 75822 151872 75828
rect 149152 74520 149204 74526
rect 149152 74462 149204 74468
rect 153212 51066 153240 155910
rect 153396 142154 153424 160126
rect 153304 142126 153424 142154
rect 153304 102134 153332 142126
rect 153292 102128 153344 102134
rect 153292 102070 153344 102076
rect 154592 75818 154620 160126
rect 154580 75812 154632 75818
rect 154580 75754 154632 75760
rect 153200 51060 153252 51066
rect 153200 51002 153252 51008
rect 155972 50998 156000 160126
rect 157340 155984 157392 155990
rect 157340 155926 157392 155932
rect 157352 77246 157380 155926
rect 157444 102066 157472 160126
rect 158088 160126 158424 160154
rect 158732 160126 159436 160154
rect 160112 160126 160448 160154
rect 158088 155990 158116 160126
rect 158076 155984 158128 155990
rect 158076 155926 158128 155932
rect 157432 102060 157484 102066
rect 157432 102002 157484 102008
rect 157340 77240 157392 77246
rect 157340 77182 157392 77188
rect 158732 52426 158760 160126
rect 160112 103494 160140 160126
rect 161480 155984 161532 155990
rect 161480 155926 161532 155932
rect 160100 103488 160152 103494
rect 160100 103430 160152 103436
rect 158720 52420 158772 52426
rect 158720 52362 158772 52368
rect 161492 52358 161520 155926
rect 161676 142154 161704 160262
rect 162136 160126 162472 160154
rect 162872 160126 163484 160154
rect 164344 160126 164496 160154
rect 165172 160126 165508 160154
rect 165632 160126 166520 160154
rect 167012 160126 167532 160154
rect 168392 160126 168636 160154
rect 169220 160126 169648 160154
rect 169772 160126 170660 160154
rect 171152 160126 171672 160154
rect 172684 160126 172744 160154
rect 162136 155990 162164 160126
rect 162124 155984 162176 155990
rect 162124 155926 162176 155932
rect 161584 142126 161704 142154
rect 161584 77178 161612 142126
rect 162872 103426 162900 160126
rect 164240 155984 164292 155990
rect 164240 155926 164292 155932
rect 162860 103420 162912 103426
rect 162860 103362 162912 103368
rect 161572 77172 161624 77178
rect 161572 77114 161624 77120
rect 164252 53786 164280 155926
rect 164344 78674 164372 160126
rect 165172 155990 165200 160126
rect 165160 155984 165212 155990
rect 165160 155926 165212 155932
rect 165632 104854 165660 160126
rect 165620 104848 165672 104854
rect 165620 104790 165672 104796
rect 167012 80034 167040 160126
rect 167000 80028 167052 80034
rect 167000 79970 167052 79976
rect 164332 78668 164384 78674
rect 164332 78610 164384 78616
rect 164240 53780 164292 53786
rect 164240 53722 164292 53728
rect 168392 53718 168420 160126
rect 169220 142154 169248 160126
rect 168484 142126 169248 142154
rect 168484 106282 168512 142126
rect 168472 106276 168524 106282
rect 168472 106218 168524 106224
rect 169772 79966 169800 160126
rect 169760 79960 169812 79966
rect 169760 79902 169812 79908
rect 171152 55214 171180 160126
rect 172520 155984 172572 155990
rect 172520 155926 172572 155932
rect 172532 81394 172560 155926
rect 172716 142154 172744 160126
rect 173360 160126 173696 160154
rect 173912 160126 174708 160154
rect 175292 160126 175720 160154
rect 176732 160126 176792 160154
rect 173360 155990 173388 160126
rect 173348 155984 173400 155990
rect 173348 155926 173400 155932
rect 172624 142126 172744 142154
rect 172624 106214 172652 142126
rect 172612 106208 172664 106214
rect 172612 106150 172664 106156
rect 172520 81388 172572 81394
rect 172520 81330 172572 81336
rect 173912 56574 173940 160126
rect 175292 107642 175320 160126
rect 176660 155984 176712 155990
rect 176660 155926 176712 155932
rect 175280 107636 175332 107642
rect 175280 107578 175332 107584
rect 173900 56568 173952 56574
rect 173900 56510 173952 56516
rect 176672 56506 176700 155926
rect 176764 81326 176792 160126
rect 177408 160126 177744 160154
rect 178052 160126 178756 160154
rect 179432 160126 179860 160154
rect 180872 160126 180932 160154
rect 177408 155990 177436 160126
rect 177396 155984 177448 155990
rect 177396 155926 177448 155932
rect 178052 107574 178080 160126
rect 178040 107568 178092 107574
rect 178040 107510 178092 107516
rect 179432 82822 179460 160126
rect 180904 155938 180932 160126
rect 180812 155910 180932 155938
rect 181088 160126 181884 160154
rect 182192 160126 182896 160154
rect 183572 160126 183908 160154
rect 184920 160126 185072 160154
rect 179420 82816 179472 82822
rect 179420 82758 179472 82764
rect 176752 81320 176804 81326
rect 176752 81262 176804 81268
rect 180812 57934 180840 155910
rect 181088 142154 181116 160126
rect 180904 142126 181116 142154
rect 180904 109002 180932 142126
rect 180892 108996 180944 109002
rect 180892 108938 180944 108944
rect 182192 82754 182220 160126
rect 182180 82748 182232 82754
rect 182180 82690 182232 82696
rect 180800 57928 180852 57934
rect 180800 57870 180852 57876
rect 183572 57866 183600 160126
rect 184940 155984 184992 155990
rect 184940 155926 184992 155932
rect 184952 84182 184980 155926
rect 185044 108934 185072 160126
rect 185596 160126 185932 160154
rect 186332 160126 186944 160154
rect 187804 160126 187956 160154
rect 188632 160126 188968 160154
rect 189092 160126 189980 160154
rect 190472 160126 190992 160154
rect 191944 160126 192096 160154
rect 192772 160126 193108 160154
rect 193232 160126 194120 160154
rect 194612 160126 195132 160154
rect 195992 160126 196144 160154
rect 196268 160126 197156 160154
rect 197372 160126 198168 160154
rect 198752 160126 199180 160154
rect 200192 160126 200252 160154
rect 185596 155990 185624 160126
rect 185584 155984 185636 155990
rect 185584 155926 185636 155932
rect 185032 108928 185084 108934
rect 185032 108870 185084 108876
rect 184940 84176 184992 84182
rect 184940 84118 184992 84124
rect 186332 59362 186360 160126
rect 187700 155984 187752 155990
rect 187700 155926 187752 155932
rect 187712 85542 187740 155926
rect 187804 110430 187832 160126
rect 188632 155990 188660 160126
rect 188620 155984 188672 155990
rect 188620 155926 188672 155932
rect 187792 110424 187844 110430
rect 187792 110366 187844 110372
rect 187700 85536 187752 85542
rect 187700 85478 187752 85484
rect 189092 60722 189120 160126
rect 190472 111790 190500 160126
rect 191840 153740 191892 153746
rect 191840 153682 191892 153688
rect 190460 111784 190512 111790
rect 190460 111726 190512 111732
rect 189080 60716 189132 60722
rect 189080 60658 189132 60664
rect 191852 60654 191880 153682
rect 191944 85474 191972 160126
rect 192772 153746 192800 160126
rect 192760 153740 192812 153746
rect 192760 153682 192812 153688
rect 193232 111722 193260 160126
rect 193220 111716 193272 111722
rect 193220 111658 193272 111664
rect 194612 86970 194640 160126
rect 194600 86964 194652 86970
rect 194600 86906 194652 86912
rect 191932 85468 191984 85474
rect 191932 85410 191984 85416
rect 195992 62082 196020 160126
rect 196268 142154 196296 160126
rect 196084 142126 196296 142154
rect 196084 113150 196112 142126
rect 196072 113144 196124 113150
rect 196072 113086 196124 113092
rect 197372 86902 197400 160126
rect 197360 86896 197412 86902
rect 197360 86838 197412 86844
rect 195980 62076 196032 62082
rect 195980 62018 196032 62024
rect 198752 62014 198780 160126
rect 200120 155984 200172 155990
rect 200120 155926 200172 155932
rect 200132 88330 200160 155926
rect 200224 113082 200252 160126
rect 200868 160126 201204 160154
rect 201512 160126 202216 160154
rect 202892 160126 203320 160154
rect 204332 160126 204392 160154
rect 200868 155990 200896 160126
rect 200856 155984 200908 155990
rect 200856 155926 200908 155932
rect 200212 113076 200264 113082
rect 200212 113018 200264 113024
rect 200120 88324 200172 88330
rect 200120 88266 200172 88272
rect 201512 63510 201540 160126
rect 202892 114510 202920 160126
rect 204260 155984 204312 155990
rect 204260 155926 204312 155932
rect 202880 114504 202932 114510
rect 202880 114446 202932 114452
rect 201500 63504 201552 63510
rect 201500 63446 201552 63452
rect 204272 63442 204300 155926
rect 204364 88262 204392 160126
rect 205008 160126 205344 160154
rect 205652 160126 206356 160154
rect 207032 160126 207368 160154
rect 208380 160126 208440 160154
rect 205008 155990 205036 160126
rect 204996 155984 205048 155990
rect 204996 155926 205048 155932
rect 205652 115938 205680 160126
rect 205640 115932 205692 115938
rect 205640 115874 205692 115880
rect 207032 89690 207060 160126
rect 207020 89684 207072 89690
rect 207020 89626 207072 89632
rect 204352 88256 204404 88262
rect 204352 88198 204404 88204
rect 208412 64870 208440 160126
rect 208504 160126 209392 160154
rect 209792 160126 210404 160154
rect 211172 160126 211416 160154
rect 211540 160126 212428 160154
rect 212552 160126 213440 160154
rect 214208 160126 214544 160154
rect 215556 160126 215892 160154
rect 208504 115870 208532 160126
rect 208492 115864 208544 115870
rect 208492 115806 208544 115812
rect 209792 91050 209820 160126
rect 209780 91044 209832 91050
rect 209780 90986 209832 90992
rect 211172 66162 211200 160126
rect 211540 142154 211568 160126
rect 211264 142126 211568 142154
rect 211264 117230 211292 142126
rect 211252 117224 211304 117230
rect 211252 117166 211304 117172
rect 212552 90982 212580 160126
rect 214208 158506 214236 160126
rect 215864 158545 215892 160126
rect 217244 160126 217580 160154
rect 219452 160126 219604 160154
rect 220616 160126 220768 160154
rect 217244 158914 217272 160126
rect 217232 158908 217284 158914
rect 217232 158850 217284 158856
rect 219452 158710 219480 160126
rect 219440 158704 219492 158710
rect 219440 158646 219492 158652
rect 215850 158536 215906 158545
rect 214196 158500 214248 158506
rect 215850 158471 215906 158480
rect 214196 158442 214248 158448
rect 220740 158409 220768 160126
rect 221292 160126 221628 160154
rect 222304 160126 222640 160154
rect 223652 160126 223712 160154
rect 221292 158438 221320 160126
rect 221280 158432 221332 158438
rect 220726 158400 220782 158409
rect 221280 158374 221332 158380
rect 220726 158335 220782 158344
rect 222304 158137 222332 160126
rect 223684 158273 223712 160126
rect 224328 160126 224664 160154
rect 225340 160126 225676 160154
rect 226780 160126 227116 160154
rect 227792 160126 228128 160154
rect 228804 160126 228956 160154
rect 229816 160126 230152 160154
rect 230828 160126 231164 160154
rect 231840 160126 231900 160154
rect 224328 158846 224356 160126
rect 224316 158840 224368 158846
rect 224316 158782 224368 158788
rect 225340 158574 225368 160126
rect 225328 158568 225380 158574
rect 225328 158510 225380 158516
rect 223670 158264 223726 158273
rect 227088 158234 227116 160126
rect 223670 158199 223726 158208
rect 227076 158228 227128 158234
rect 227076 158170 227128 158176
rect 222290 158128 222346 158137
rect 222290 158063 222346 158072
rect 228100 157962 228128 160126
rect 228928 158137 228956 160126
rect 230124 158302 230152 160126
rect 231136 158438 231164 160126
rect 231124 158432 231176 158438
rect 231124 158374 231176 158380
rect 230112 158296 230164 158302
rect 230112 158238 230164 158244
rect 228914 158128 228970 158137
rect 228914 158063 228970 158072
rect 228088 157956 228140 157962
rect 228088 157898 228140 157904
rect 231872 157826 231900 160126
rect 232516 160126 232852 160154
rect 233528 160126 233864 160154
rect 234632 160126 234876 160154
rect 235888 160126 235948 160154
rect 232516 157894 232544 160126
rect 233528 159254 233556 160126
rect 233516 159248 233568 159254
rect 233516 159190 233568 159196
rect 234632 158166 234660 160126
rect 235920 158710 235948 160126
rect 236564 160126 236900 160154
rect 237668 160126 238004 160154
rect 239016 160126 239352 160154
rect 240028 160126 240088 160154
rect 235908 158704 235960 158710
rect 235908 158646 235960 158652
rect 234620 158160 234672 158166
rect 234620 158102 234672 158108
rect 236564 158098 236592 160126
rect 236552 158092 236604 158098
rect 236552 158034 236604 158040
rect 237668 158030 237696 160126
rect 239324 158574 239352 160126
rect 240060 158846 240088 160126
rect 240704 160126 241040 160154
rect 242052 160126 242388 160154
rect 243064 160126 243400 160154
rect 240704 159322 240732 160126
rect 240692 159316 240744 159322
rect 240692 159258 240744 159264
rect 240048 158840 240100 158846
rect 240048 158782 240100 158788
rect 239312 158568 239364 158574
rect 239312 158510 239364 158516
rect 242360 158506 242388 160126
rect 242808 159452 242860 159458
rect 242808 159394 242860 159400
rect 242348 158500 242400 158506
rect 242348 158442 242400 158448
rect 242820 158438 242848 159394
rect 243372 158914 243400 160126
rect 243740 160126 244076 160154
rect 245088 160126 245424 160154
rect 246100 160126 246436 160154
rect 247112 160126 247172 160154
rect 248124 160126 248276 160154
rect 249228 160126 249564 160154
rect 243740 159186 243768 160126
rect 244280 159384 244332 159390
rect 244280 159326 244332 159332
rect 243728 159180 243780 159186
rect 243728 159122 243780 159128
rect 243360 158908 243412 158914
rect 243360 158850 243412 158856
rect 244292 158710 244320 159326
rect 244280 158704 244332 158710
rect 244280 158646 244332 158652
rect 245396 158438 245424 160126
rect 246408 159186 246436 160126
rect 246396 159180 246448 159186
rect 246396 159122 246448 159128
rect 247144 158982 247172 160126
rect 247132 158976 247184 158982
rect 247132 158918 247184 158924
rect 248248 158710 248276 160126
rect 249536 158982 249564 160126
rect 249904 160126 250240 160154
rect 251252 160126 251312 160154
rect 249904 159118 249932 160126
rect 249892 159112 249944 159118
rect 249892 159054 249944 159060
rect 249524 158976 249576 158982
rect 249524 158918 249576 158924
rect 248236 158704 248288 158710
rect 248236 158646 248288 158652
rect 251284 158642 251312 160126
rect 251928 160126 252264 160154
rect 253276 160126 253612 160154
rect 251272 158636 251324 158642
rect 251272 158578 251324 158584
rect 242808 158432 242860 158438
rect 242808 158374 242860 158380
rect 245384 158432 245436 158438
rect 245384 158374 245436 158380
rect 237656 158024 237708 158030
rect 251928 158001 251956 160126
rect 253584 159118 253612 160126
rect 253952 160126 254288 160154
rect 255300 160126 255636 160154
rect 256312 160126 256648 160154
rect 253572 159112 253624 159118
rect 253572 159054 253624 159060
rect 253952 159050 253980 160126
rect 253940 159044 253992 159050
rect 253940 158986 253992 158992
rect 255608 158642 255636 160126
rect 256620 159254 256648 160126
rect 256988 160126 257324 160154
rect 258184 160126 258336 160154
rect 259348 160126 259408 160154
rect 256608 159248 256660 159254
rect 256608 159190 256660 159196
rect 255596 158636 255648 158642
rect 255596 158578 255648 158584
rect 256988 158370 257016 160126
rect 256976 158364 257028 158370
rect 256976 158306 257028 158312
rect 258184 158273 258212 160126
rect 259380 159050 259408 160126
rect 260380 160132 260432 160138
rect 260380 160074 260432 160080
rect 259368 159044 259420 159050
rect 259368 158986 259420 158992
rect 258170 158264 258226 158273
rect 260392 158234 260420 160074
rect 263612 158846 263640 297871
rect 263704 160138 263732 298007
rect 264336 297968 264388 297974
rect 264336 297910 264388 297916
rect 264244 296744 264296 296750
rect 264244 296686 264296 296692
rect 263692 160132 263744 160138
rect 263692 160074 263744 160080
rect 263600 158840 263652 158846
rect 263600 158782 263652 158788
rect 258170 158199 258226 158208
rect 260380 158228 260432 158234
rect 260380 158170 260432 158176
rect 237656 157966 237708 157972
rect 251914 157992 251970 158001
rect 264256 157962 264284 296686
rect 264348 189990 264376 297910
rect 265084 235346 265112 298007
rect 265360 297974 265388 298007
rect 265348 297968 265400 297974
rect 265348 297910 265400 297916
rect 265072 235340 265124 235346
rect 265072 235282 265124 235288
rect 264336 189984 264388 189990
rect 264336 189926 264388 189932
rect 266372 158914 266400 298007
rect 266450 297936 266506 297945
rect 266450 297871 266506 297880
rect 266464 159186 266492 297871
rect 267844 235278 267872 298007
rect 268014 297936 268070 297945
rect 268014 297871 268070 297880
rect 268028 296750 268056 297871
rect 269776 297022 269804 298007
rect 269764 297016 269816 297022
rect 269764 296958 269816 296964
rect 268016 296744 268068 296750
rect 268016 296686 268068 296692
rect 267832 235272 267884 235278
rect 267832 235214 267884 235220
rect 266452 159180 266504 159186
rect 266452 159122 266504 159128
rect 266360 158908 266412 158914
rect 266360 158850 266412 158856
rect 270512 158302 270540 298007
rect 270590 297936 270646 297945
rect 270590 297871 270646 297880
rect 270604 158982 270632 297871
rect 271892 236774 271920 298007
rect 271880 236768 271932 236774
rect 271880 236710 271932 236716
rect 273272 159118 273300 298007
rect 273350 297936 273406 297945
rect 273350 297871 273406 297880
rect 273364 159458 273392 297871
rect 273442 297800 273498 297809
rect 273442 297735 273498 297744
rect 273456 236842 273484 297735
rect 273444 236836 273496 236842
rect 273444 236778 273496 236784
rect 273352 159452 273404 159458
rect 273352 159394 273404 159400
rect 274652 159254 274680 298007
rect 275284 297968 275336 297974
rect 275284 297910 275336 297916
rect 275296 232626 275324 297910
rect 276032 297226 276060 298007
rect 276768 297974 276796 298007
rect 276756 297968 276808 297974
rect 276756 297910 276808 297916
rect 276020 297220 276072 297226
rect 276020 297162 276072 297168
rect 276662 296984 276718 296993
rect 276662 296919 276718 296928
rect 275284 232620 275336 232626
rect 275284 232562 275336 232568
rect 276676 224942 276704 296919
rect 276664 224936 276716 224942
rect 276664 224878 276716 224884
rect 277504 204270 277532 298007
rect 277492 204264 277544 204270
rect 277492 204206 277544 204212
rect 274640 159248 274692 159254
rect 274640 159190 274692 159196
rect 273260 159112 273312 159118
rect 273260 159054 273312 159060
rect 278792 159050 278820 298007
rect 280172 240990 280200 298007
rect 282184 297968 282236 297974
rect 282184 297910 282236 297916
rect 280160 240984 280212 240990
rect 280160 240926 280212 240932
rect 282196 232898 282224 297910
rect 282184 232892 282236 232898
rect 282184 232834 282236 232840
rect 282932 159390 282960 298007
rect 285968 297974 285996 298007
rect 285956 297968 286008 297974
rect 285956 297910 286008 297916
rect 286324 296812 286376 296818
rect 286324 296754 286376 296760
rect 284944 296744 284996 296750
rect 284944 296686 284996 296692
rect 284956 232966 284984 296686
rect 284944 232960 284996 232966
rect 284944 232902 284996 232908
rect 282920 159384 282972 159390
rect 282920 159326 282972 159332
rect 278780 159044 278832 159050
rect 278780 158986 278832 158992
rect 270592 158976 270644 158982
rect 270592 158918 270644 158924
rect 286336 158574 286364 296754
rect 287624 296750 287652 298007
rect 287704 297968 287756 297974
rect 287704 297910 287756 297916
rect 287612 296744 287664 296750
rect 287612 296686 287664 296692
rect 286324 158568 286376 158574
rect 286324 158510 286376 158516
rect 287716 158506 287744 297910
rect 289084 296948 289136 296954
rect 289084 296890 289136 296896
rect 287704 158500 287756 158506
rect 287704 158442 287756 158448
rect 289096 158438 289124 296890
rect 290016 296818 290044 298007
rect 290004 296812 290056 296818
rect 290004 296754 290056 296760
rect 291844 296812 291896 296818
rect 291844 296754 291896 296760
rect 291856 211138 291884 296754
rect 292592 240922 292620 298007
rect 295352 297974 295380 298007
rect 295340 297968 295392 297974
rect 295340 297910 295392 297916
rect 294604 297016 294656 297022
rect 294604 296958 294656 296964
rect 292580 240916 292632 240922
rect 292580 240858 292632 240864
rect 294616 213926 294644 296958
rect 298480 296954 298508 298007
rect 298468 296948 298520 296954
rect 298468 296890 298520 296896
rect 300124 296948 300176 296954
rect 300124 296890 300176 296896
rect 295984 296880 296036 296886
rect 295984 296822 296036 296828
rect 294604 213920 294656 213926
rect 294604 213862 294656 213868
rect 291844 211132 291896 211138
rect 291844 211074 291896 211080
rect 295996 158710 296024 296822
rect 298744 296744 298796 296750
rect 298744 296686 298796 296692
rect 298756 216646 298784 296686
rect 300136 218006 300164 296890
rect 300872 296818 300900 298007
rect 302344 297022 302372 298007
rect 302884 297084 302936 297090
rect 302884 297026 302936 297032
rect 302332 297016 302384 297022
rect 302332 296958 302384 296964
rect 300860 296812 300912 296818
rect 300860 296754 300912 296760
rect 300124 218000 300176 218006
rect 300124 217942 300176 217948
rect 298744 216640 298796 216646
rect 298744 216582 298796 216588
rect 295984 158704 296036 158710
rect 295984 158646 296036 158652
rect 302896 158642 302924 297026
rect 305104 296886 305132 298007
rect 305644 297016 305696 297022
rect 305644 296958 305696 296964
rect 305092 296880 305144 296886
rect 305092 296822 305144 296828
rect 304264 296812 304316 296818
rect 304264 296754 304316 296760
rect 304276 232558 304304 296754
rect 304264 232552 304316 232558
rect 304264 232494 304316 232500
rect 305656 223582 305684 296958
rect 308600 296750 308628 298007
rect 310992 296954 311020 298007
rect 310980 296948 311032 296954
rect 310980 296890 311032 296896
rect 308588 296744 308640 296750
rect 308588 296686 308640 296692
rect 313292 240786 313320 298007
rect 315776 297090 315804 298007
rect 315764 297084 315816 297090
rect 315764 297026 315816 297032
rect 317432 296818 317460 298007
rect 320928 297022 320956 298007
rect 320916 297016 320968 297022
rect 320916 296958 320968 296964
rect 317420 296812 317472 296818
rect 317420 296754 317472 296760
rect 313280 240780 313332 240786
rect 313280 240722 313332 240728
rect 322952 231266 322980 298007
rect 322940 231260 322992 231266
rect 322940 231202 322992 231208
rect 325712 231130 325740 298007
rect 343232 298007 343234 298016
rect 343362 298072 343364 298081
rect 343416 298072 343418 298081
rect 343362 298007 343418 298016
rect 343180 297978 343232 297984
rect 325700 231124 325752 231130
rect 325700 231066 325752 231072
rect 305644 223576 305696 223582
rect 305644 223518 305696 223524
rect 302884 158636 302936 158642
rect 302884 158578 302936 158584
rect 289084 158432 289136 158438
rect 289084 158374 289136 158380
rect 270500 158296 270552 158302
rect 270500 158238 270552 158244
rect 251914 157927 251970 157936
rect 264244 157956 264296 157962
rect 264244 157898 264296 157904
rect 232504 157888 232556 157894
rect 232504 157830 232556 157836
rect 231860 157820 231912 157826
rect 231860 157762 231912 157768
rect 256700 120080 256752 120086
rect 256700 120022 256752 120028
rect 342260 120080 342312 120086
rect 342260 120022 342312 120028
rect 256712 119513 256740 120022
rect 342272 119513 342300 120022
rect 256698 119504 256754 119513
rect 256698 119439 256754 119448
rect 342258 119504 342314 119513
rect 342258 119439 342314 119448
rect 256698 118688 256754 118697
rect 256698 118623 256700 118632
rect 256752 118623 256754 118632
rect 342258 118688 342314 118697
rect 342258 118623 342314 118632
rect 342352 118652 342404 118658
rect 256700 118594 256752 118600
rect 342272 118590 342300 118623
rect 342352 118594 342404 118600
rect 256792 118584 256844 118590
rect 256792 118526 256844 118532
rect 342260 118584 342312 118590
rect 342260 118526 342312 118532
rect 256804 117881 256832 118526
rect 342364 117881 342392 118594
rect 256790 117872 256846 117881
rect 256790 117807 256846 117816
rect 342350 117872 342406 117881
rect 342350 117807 342406 117816
rect 256700 117292 256752 117298
rect 256700 117234 256752 117240
rect 342352 117292 342404 117298
rect 342352 117234 342404 117240
rect 256712 117065 256740 117234
rect 256792 117224 256844 117230
rect 256792 117166 256844 117172
rect 342260 117224 342312 117230
rect 342260 117166 342312 117172
rect 256698 117056 256754 117065
rect 256698 116991 256754 117000
rect 256804 116249 256832 117166
rect 342272 117065 342300 117166
rect 342258 117056 342314 117065
rect 342258 116991 342314 117000
rect 342364 116249 342392 117234
rect 256790 116240 256846 116249
rect 256790 116175 256846 116184
rect 342350 116240 342406 116249
rect 342350 116175 342406 116184
rect 256792 115932 256844 115938
rect 256792 115874 256844 115880
rect 342260 115932 342312 115938
rect 342260 115874 342312 115880
rect 256700 115864 256752 115870
rect 256700 115806 256752 115812
rect 256712 115433 256740 115806
rect 256698 115424 256754 115433
rect 256698 115359 256754 115368
rect 256804 114617 256832 115874
rect 342272 115433 342300 115874
rect 342352 115864 342404 115870
rect 342352 115806 342404 115812
rect 342258 115424 342314 115433
rect 342258 115359 342314 115368
rect 342364 114617 342392 115806
rect 256790 114608 256846 114617
rect 256790 114543 256846 114552
rect 342350 114608 342406 114617
rect 342350 114543 342406 114552
rect 256700 114504 256752 114510
rect 256700 114446 256752 114452
rect 342260 114504 342312 114510
rect 342260 114446 342312 114452
rect 256712 113801 256740 114446
rect 342272 113801 342300 114446
rect 256698 113792 256754 113801
rect 256698 113727 256754 113736
rect 342258 113792 342314 113801
rect 342258 113727 342314 113736
rect 256792 113144 256844 113150
rect 256698 113112 256754 113121
rect 342260 113144 342312 113150
rect 256792 113086 256844 113092
rect 342258 113112 342260 113121
rect 342312 113112 342314 113121
rect 256698 113047 256700 113056
rect 256752 113047 256754 113056
rect 256700 113018 256752 113024
rect 256804 112305 256832 113086
rect 342258 113047 342314 113056
rect 342352 113076 342404 113082
rect 342352 113018 342404 113024
rect 342364 112305 342392 113018
rect 256790 112296 256846 112305
rect 256790 112231 256846 112240
rect 342350 112296 342406 112305
rect 342350 112231 342406 112240
rect 256792 111784 256844 111790
rect 256792 111726 256844 111732
rect 342260 111784 342312 111790
rect 342260 111726 342312 111732
rect 256700 111716 256752 111722
rect 256700 111658 256752 111664
rect 256712 111489 256740 111658
rect 256698 111480 256754 111489
rect 256698 111415 256754 111424
rect 256804 110673 256832 111726
rect 342272 111489 342300 111726
rect 342352 111716 342404 111722
rect 342352 111658 342404 111664
rect 342258 111480 342314 111489
rect 342258 111415 342314 111424
rect 342364 110673 342392 111658
rect 256790 110664 256846 110673
rect 256790 110599 256846 110608
rect 342350 110664 342406 110673
rect 342350 110599 342406 110608
rect 256700 110424 256752 110430
rect 256700 110366 256752 110372
rect 342260 110424 342312 110430
rect 342260 110366 342312 110372
rect 256712 109857 256740 110366
rect 342272 109857 342300 110366
rect 256698 109848 256754 109857
rect 256698 109783 256754 109792
rect 342258 109848 342314 109857
rect 342258 109783 342314 109792
rect 256698 109032 256754 109041
rect 342258 109032 342314 109041
rect 256698 108967 256754 108976
rect 256792 108996 256844 109002
rect 256712 108934 256740 108967
rect 342258 108967 342260 108976
rect 256792 108938 256844 108944
rect 342312 108967 342314 108976
rect 342260 108938 342312 108944
rect 256700 108928 256752 108934
rect 256700 108870 256752 108876
rect 256804 108225 256832 108938
rect 342352 108928 342404 108934
rect 342352 108870 342404 108876
rect 342364 108225 342392 108870
rect 256790 108216 256846 108225
rect 256790 108151 256846 108160
rect 342350 108216 342406 108225
rect 342350 108151 342406 108160
rect 256792 107636 256844 107642
rect 256792 107578 256844 107584
rect 342260 107636 342312 107642
rect 342260 107578 342312 107584
rect 256700 107568 256752 107574
rect 256700 107510 256752 107516
rect 256712 107409 256740 107510
rect 256698 107400 256754 107409
rect 256698 107335 256754 107344
rect 256804 106729 256832 107578
rect 342272 107409 342300 107578
rect 342352 107568 342404 107574
rect 342352 107510 342404 107516
rect 342258 107400 342314 107409
rect 342258 107335 342314 107344
rect 342364 106729 342392 107510
rect 256790 106720 256846 106729
rect 256790 106655 256846 106664
rect 342350 106720 342406 106729
rect 342350 106655 342406 106664
rect 256792 106276 256844 106282
rect 256792 106218 256844 106224
rect 342352 106276 342404 106282
rect 342352 106218 342404 106224
rect 256700 106208 256752 106214
rect 256700 106150 256752 106156
rect 256712 105913 256740 106150
rect 256698 105904 256754 105913
rect 256698 105839 256754 105848
rect 256804 105097 256832 106218
rect 342260 106208 342312 106214
rect 342260 106150 342312 106156
rect 342272 105913 342300 106150
rect 342258 105904 342314 105913
rect 342258 105839 342314 105848
rect 342364 105097 342392 106218
rect 256790 105088 256846 105097
rect 256790 105023 256846 105032
rect 342350 105088 342406 105097
rect 342350 105023 342406 105032
rect 256700 104848 256752 104854
rect 256700 104790 256752 104796
rect 342260 104848 342312 104854
rect 342260 104790 342312 104796
rect 256712 104281 256740 104790
rect 342272 104281 342300 104790
rect 256698 104272 256754 104281
rect 256698 104207 256754 104216
rect 342258 104272 342314 104281
rect 342258 104207 342314 104216
rect 256792 103488 256844 103494
rect 256698 103456 256754 103465
rect 342260 103488 342312 103494
rect 256792 103430 256844 103436
rect 342258 103456 342260 103465
rect 342312 103456 342314 103465
rect 256698 103391 256700 103400
rect 256752 103391 256754 103400
rect 256700 103362 256752 103368
rect 256804 102649 256832 103430
rect 342258 103391 342314 103400
rect 342352 103420 342404 103426
rect 342352 103362 342404 103368
rect 342364 102649 342392 103362
rect 256790 102640 256846 102649
rect 256790 102575 256846 102584
rect 342350 102640 342406 102649
rect 342350 102575 342406 102584
rect 256792 102128 256844 102134
rect 256792 102070 256844 102076
rect 342260 102128 342312 102134
rect 342260 102070 342312 102076
rect 256700 102060 256752 102066
rect 256700 102002 256752 102008
rect 256712 101833 256740 102002
rect 256698 101824 256754 101833
rect 256698 101759 256754 101768
rect 256804 101017 256832 102070
rect 342272 101833 342300 102070
rect 342352 102060 342404 102066
rect 342352 102002 342404 102008
rect 342258 101824 342314 101833
rect 342258 101759 342314 101768
rect 342364 101017 342392 102002
rect 256790 101008 256846 101017
rect 256790 100943 256846 100952
rect 342350 101008 342406 101017
rect 342350 100943 342406 100952
rect 256792 100700 256844 100706
rect 256792 100642 256844 100648
rect 342260 100700 342312 100706
rect 342260 100642 342312 100648
rect 256700 100632 256752 100638
rect 256700 100574 256752 100580
rect 256712 100337 256740 100574
rect 256698 100328 256754 100337
rect 256698 100263 256754 100272
rect 256804 99521 256832 100642
rect 342272 100337 342300 100642
rect 342352 100632 342404 100638
rect 342352 100574 342404 100580
rect 342258 100328 342314 100337
rect 342258 100263 342314 100272
rect 342364 99521 342392 100574
rect 256790 99512 256846 99521
rect 256790 99447 256846 99456
rect 342350 99512 342406 99521
rect 342350 99447 342406 99456
rect 256700 99340 256752 99346
rect 256700 99282 256752 99288
rect 342260 99340 342312 99346
rect 342260 99282 342312 99288
rect 256712 98705 256740 99282
rect 342272 98705 342300 99282
rect 256698 98696 256754 98705
rect 256698 98631 256754 98640
rect 342258 98696 342314 98705
rect 342258 98631 342314 98640
rect 256792 97980 256844 97986
rect 256792 97922 256844 97928
rect 342260 97980 342312 97986
rect 342260 97922 342312 97928
rect 256700 97912 256752 97918
rect 256698 97880 256700 97889
rect 256752 97880 256754 97889
rect 256698 97815 256754 97824
rect 256804 97073 256832 97922
rect 342272 97889 342300 97922
rect 342352 97912 342404 97918
rect 342258 97880 342314 97889
rect 342352 97854 342404 97860
rect 342258 97815 342314 97824
rect 342364 97073 342392 97854
rect 256790 97064 256846 97073
rect 256790 96999 256846 97008
rect 342350 97064 342406 97073
rect 342350 96999 342406 97008
rect 256792 96620 256844 96626
rect 256792 96562 256844 96568
rect 342260 96620 342312 96626
rect 342260 96562 342312 96568
rect 256700 96552 256752 96558
rect 256700 96494 256752 96500
rect 256712 96257 256740 96494
rect 256698 96248 256754 96257
rect 256698 96183 256754 96192
rect 256804 95441 256832 96562
rect 342272 96257 342300 96562
rect 342352 96552 342404 96558
rect 342352 96494 342404 96500
rect 342258 96248 342314 96257
rect 342258 96183 342314 96192
rect 342364 95441 342392 96494
rect 256790 95432 256846 95441
rect 256790 95367 256846 95376
rect 342350 95432 342406 95441
rect 342350 95367 342406 95376
rect 256700 95192 256752 95198
rect 256700 95134 256752 95140
rect 342260 95192 342312 95198
rect 342260 95134 342312 95140
rect 256712 94625 256740 95134
rect 342272 94625 342300 95134
rect 256698 94616 256754 94625
rect 256698 94551 256754 94560
rect 342258 94616 342314 94625
rect 342258 94551 342314 94560
rect 256792 93832 256844 93838
rect 256698 93800 256754 93809
rect 342260 93832 342312 93838
rect 256792 93774 256844 93780
rect 342258 93800 342260 93809
rect 342312 93800 342314 93809
rect 256698 93735 256700 93744
rect 256752 93735 256754 93744
rect 256700 93706 256752 93712
rect 256804 93129 256832 93774
rect 342258 93735 342314 93744
rect 342352 93764 342404 93770
rect 342352 93706 342404 93712
rect 342364 93129 342392 93706
rect 256790 93120 256846 93129
rect 256790 93055 256846 93064
rect 342350 93120 342406 93129
rect 342350 93055 342406 93064
rect 256792 92472 256844 92478
rect 256792 92414 256844 92420
rect 342260 92472 342312 92478
rect 342260 92414 342312 92420
rect 256700 92404 256752 92410
rect 256700 92346 256752 92352
rect 256712 92313 256740 92346
rect 256698 92304 256754 92313
rect 256698 92239 256754 92248
rect 256804 91497 256832 92414
rect 342272 92313 342300 92414
rect 342352 92404 342404 92410
rect 342352 92346 342404 92352
rect 342258 92304 342314 92313
rect 342258 92239 342314 92248
rect 342364 91497 342392 92346
rect 256790 91488 256846 91497
rect 256790 91423 256846 91432
rect 342350 91488 342406 91497
rect 342350 91423 342406 91432
rect 256792 91044 256844 91050
rect 256792 90986 256844 90992
rect 342260 91044 342312 91050
rect 342260 90986 342312 90992
rect 212540 90976 212592 90982
rect 212540 90918 212592 90924
rect 256700 90976 256752 90982
rect 256700 90918 256752 90924
rect 256712 90681 256740 90918
rect 256698 90672 256754 90681
rect 256698 90607 256754 90616
rect 256804 89865 256832 90986
rect 342272 90681 342300 90986
rect 342352 90976 342404 90982
rect 342352 90918 342404 90924
rect 342258 90672 342314 90681
rect 342258 90607 342314 90616
rect 342364 89865 342392 90918
rect 256790 89856 256846 89865
rect 256790 89791 256846 89800
rect 342350 89856 342406 89865
rect 342350 89791 342406 89800
rect 256700 89684 256752 89690
rect 256700 89626 256752 89632
rect 342260 89684 342312 89690
rect 342260 89626 342312 89632
rect 256712 89049 256740 89626
rect 342272 89049 342300 89626
rect 256698 89040 256754 89049
rect 256698 88975 256754 88984
rect 342258 89040 342314 89049
rect 342258 88975 342314 88984
rect 256792 88324 256844 88330
rect 256792 88266 256844 88272
rect 342260 88324 342312 88330
rect 342260 88266 342312 88272
rect 256700 88256 256752 88262
rect 256698 88224 256700 88233
rect 256752 88224 256754 88233
rect 256698 88159 256754 88168
rect 256804 87417 256832 88266
rect 342272 88233 342300 88266
rect 342352 88256 342404 88262
rect 342258 88224 342314 88233
rect 342352 88198 342404 88204
rect 342258 88159 342314 88168
rect 342364 87417 342392 88198
rect 256790 87408 256846 87417
rect 256790 87343 256846 87352
rect 342350 87408 342406 87417
rect 342350 87343 342406 87352
rect 256792 86964 256844 86970
rect 256792 86906 256844 86912
rect 342260 86964 342312 86970
rect 342260 86906 342312 86912
rect 256700 86896 256752 86902
rect 256700 86838 256752 86844
rect 256712 86737 256740 86838
rect 256698 86728 256754 86737
rect 256698 86663 256754 86672
rect 256804 85921 256832 86906
rect 342272 86737 342300 86906
rect 342352 86896 342404 86902
rect 342352 86838 342404 86844
rect 342258 86728 342314 86737
rect 342258 86663 342314 86672
rect 342364 85921 342392 86838
rect 256790 85912 256846 85921
rect 256790 85847 256846 85856
rect 342350 85912 342406 85921
rect 342350 85847 342406 85856
rect 256792 85536 256844 85542
rect 256792 85478 256844 85484
rect 342352 85536 342404 85542
rect 342352 85478 342404 85484
rect 256700 85468 256752 85474
rect 256700 85410 256752 85416
rect 256712 85105 256740 85410
rect 256698 85096 256754 85105
rect 256698 85031 256754 85040
rect 256804 84289 256832 85478
rect 342260 85468 342312 85474
rect 342260 85410 342312 85416
rect 342272 85105 342300 85410
rect 342258 85096 342314 85105
rect 342258 85031 342314 85040
rect 342364 84289 342392 85478
rect 256790 84280 256846 84289
rect 256790 84215 256846 84224
rect 342350 84280 342406 84289
rect 342350 84215 342406 84224
rect 256700 84176 256752 84182
rect 256700 84118 256752 84124
rect 342260 84176 342312 84182
rect 342260 84118 342312 84124
rect 256712 83473 256740 84118
rect 342272 83473 342300 84118
rect 256698 83464 256754 83473
rect 256698 83399 256754 83408
rect 342258 83464 342314 83473
rect 342258 83399 342314 83408
rect 256792 82816 256844 82822
rect 256792 82758 256844 82764
rect 342260 82816 342312 82822
rect 342260 82758 342312 82764
rect 256700 82748 256752 82754
rect 256700 82690 256752 82696
rect 256712 82657 256740 82690
rect 256698 82648 256754 82657
rect 256698 82583 256754 82592
rect 256804 81841 256832 82758
rect 342272 82657 342300 82758
rect 342352 82748 342404 82754
rect 342352 82690 342404 82696
rect 342258 82648 342314 82657
rect 342258 82583 342314 82592
rect 342364 81841 342392 82690
rect 256790 81832 256846 81841
rect 256790 81767 256846 81776
rect 342350 81832 342406 81841
rect 342350 81767 342406 81776
rect 256792 81388 256844 81394
rect 256792 81330 256844 81336
rect 342260 81388 342312 81394
rect 342260 81330 342312 81336
rect 256700 81320 256752 81326
rect 256700 81262 256752 81268
rect 256712 81025 256740 81262
rect 256698 81016 256754 81025
rect 256698 80951 256754 80960
rect 256804 80345 256832 81330
rect 342272 81025 342300 81330
rect 342352 81320 342404 81326
rect 342352 81262 342404 81268
rect 342258 81016 342314 81025
rect 342258 80951 342314 80960
rect 342364 80345 342392 81262
rect 256790 80336 256846 80345
rect 256790 80271 256846 80280
rect 342350 80336 342406 80345
rect 342350 80271 342406 80280
rect 256792 80028 256844 80034
rect 256792 79970 256844 79976
rect 342260 80028 342312 80034
rect 342260 79970 342312 79976
rect 256700 79960 256752 79966
rect 256700 79902 256752 79908
rect 256712 79529 256740 79902
rect 256698 79520 256754 79529
rect 256698 79455 256754 79464
rect 256804 78713 256832 79970
rect 342272 79529 342300 79970
rect 342352 79960 342404 79966
rect 342352 79902 342404 79908
rect 342258 79520 342314 79529
rect 342258 79455 342314 79464
rect 342364 78713 342392 79902
rect 256790 78704 256846 78713
rect 256700 78668 256752 78674
rect 342350 78704 342406 78713
rect 256790 78639 256846 78648
rect 342260 78668 342312 78674
rect 256700 78610 256752 78616
rect 342350 78639 342406 78648
rect 342260 78610 342312 78616
rect 256712 77897 256740 78610
rect 342272 77897 342300 78610
rect 256698 77888 256754 77897
rect 256698 77823 256754 77832
rect 342258 77888 342314 77897
rect 342258 77823 342314 77832
rect 256792 77240 256844 77246
rect 256792 77182 256844 77188
rect 342260 77240 342312 77246
rect 342260 77182 342312 77188
rect 256700 77172 256752 77178
rect 256700 77114 256752 77120
rect 256712 77081 256740 77114
rect 256698 77072 256754 77081
rect 256698 77007 256754 77016
rect 256804 76265 256832 77182
rect 342272 77081 342300 77182
rect 342352 77172 342404 77178
rect 342352 77114 342404 77120
rect 342258 77072 342314 77081
rect 342258 77007 342314 77016
rect 342364 76265 342392 77114
rect 256790 76256 256846 76265
rect 256790 76191 256846 76200
rect 342350 76256 342406 76265
rect 342350 76191 342406 76200
rect 256792 75880 256844 75886
rect 256792 75822 256844 75828
rect 342260 75880 342312 75886
rect 342260 75822 342312 75828
rect 256700 75812 256752 75818
rect 256700 75754 256752 75760
rect 256712 75449 256740 75754
rect 256698 75440 256754 75449
rect 256698 75375 256754 75384
rect 256804 74633 256832 75822
rect 342272 75449 342300 75822
rect 342352 75812 342404 75818
rect 342352 75754 342404 75760
rect 342258 75440 342314 75449
rect 342258 75375 342314 75384
rect 342364 74633 342392 75754
rect 256790 74624 256846 74633
rect 256790 74559 256846 74568
rect 342350 74624 342406 74633
rect 342350 74559 342406 74568
rect 256700 74520 256752 74526
rect 256700 74462 256752 74468
rect 342260 74520 342312 74526
rect 342260 74462 342312 74468
rect 256712 73817 256740 74462
rect 342272 73817 342300 74462
rect 256698 73808 256754 73817
rect 256698 73743 256754 73752
rect 342258 73808 342314 73817
rect 342258 73743 342314 73752
rect 256792 73160 256844 73166
rect 256698 73128 256754 73137
rect 342260 73160 342312 73166
rect 256792 73102 256844 73108
rect 342258 73128 342260 73137
rect 342312 73128 342314 73137
rect 256698 73063 256700 73072
rect 256752 73063 256754 73072
rect 256700 73034 256752 73040
rect 256804 72321 256832 73102
rect 342258 73063 342314 73072
rect 342352 73092 342404 73098
rect 342352 73034 342404 73040
rect 342364 72321 342392 73034
rect 256790 72312 256846 72321
rect 256790 72247 256846 72256
rect 342350 72312 342406 72321
rect 342350 72247 342406 72256
rect 256792 71732 256844 71738
rect 256792 71674 256844 71680
rect 342352 71732 342404 71738
rect 342352 71674 342404 71680
rect 256700 71664 256752 71670
rect 256700 71606 256752 71612
rect 256712 71505 256740 71606
rect 256698 71496 256754 71505
rect 256698 71431 256754 71440
rect 256804 70689 256832 71674
rect 342260 71664 342312 71670
rect 342260 71606 342312 71612
rect 342272 71505 342300 71606
rect 342258 71496 342314 71505
rect 342258 71431 342314 71440
rect 342364 70689 342392 71674
rect 256790 70680 256846 70689
rect 256790 70615 256846 70624
rect 342350 70680 342406 70689
rect 342350 70615 342406 70624
rect 256792 70372 256844 70378
rect 256792 70314 256844 70320
rect 342260 70372 342312 70378
rect 342260 70314 342312 70320
rect 256700 70304 256752 70310
rect 256700 70246 256752 70252
rect 256712 69873 256740 70246
rect 256698 69864 256754 69873
rect 256698 69799 256754 69808
rect 256804 69057 256832 70314
rect 342272 69873 342300 70314
rect 342352 70304 342404 70310
rect 342352 70246 342404 70252
rect 342258 69864 342314 69873
rect 342258 69799 342314 69808
rect 342364 69057 342392 70246
rect 256790 69048 256846 69057
rect 256700 69012 256752 69018
rect 342350 69048 342406 69057
rect 256790 68983 256846 68992
rect 342260 69012 342312 69018
rect 256700 68954 256752 68960
rect 342350 68983 342406 68992
rect 342260 68954 342312 68960
rect 256712 68241 256740 68954
rect 342272 68241 342300 68954
rect 256698 68232 256754 68241
rect 256698 68167 256754 68176
rect 342258 68232 342314 68241
rect 342258 68167 342314 68176
rect 256792 67584 256844 67590
rect 256792 67526 256844 67532
rect 342260 67584 342312 67590
rect 342260 67526 342312 67532
rect 256700 67516 256752 67522
rect 256700 67458 256752 67464
rect 256712 67425 256740 67458
rect 256698 67416 256754 67425
rect 256698 67351 256754 67360
rect 256804 66745 256832 67526
rect 342272 67425 342300 67526
rect 342352 67516 342404 67522
rect 342352 67458 342404 67464
rect 342258 67416 342314 67425
rect 342258 67351 342314 67360
rect 342364 66745 342392 67458
rect 256790 66736 256846 66745
rect 256790 66671 256846 66680
rect 342350 66736 342406 66745
rect 342350 66671 342406 66680
rect 256700 66224 256752 66230
rect 256700 66166 256752 66172
rect 342352 66224 342404 66230
rect 342352 66166 342404 66172
rect 211160 66156 211212 66162
rect 211160 66098 211212 66104
rect 256712 65929 256740 66166
rect 256792 66156 256844 66162
rect 256792 66098 256844 66104
rect 342260 66156 342312 66162
rect 342260 66098 342312 66104
rect 256698 65920 256754 65929
rect 256698 65855 256754 65864
rect 256804 65113 256832 66098
rect 342272 65929 342300 66098
rect 342258 65920 342314 65929
rect 342258 65855 342314 65864
rect 342364 65113 342392 66166
rect 256790 65104 256846 65113
rect 256790 65039 256846 65048
rect 342350 65104 342406 65113
rect 342350 65039 342406 65048
rect 208400 64864 208452 64870
rect 208400 64806 208452 64812
rect 256700 64864 256752 64870
rect 256700 64806 256752 64812
rect 342260 64864 342312 64870
rect 342260 64806 342312 64812
rect 256712 64297 256740 64806
rect 342272 64297 342300 64806
rect 256698 64288 256754 64297
rect 256698 64223 256754 64232
rect 342258 64288 342314 64297
rect 342258 64223 342314 64232
rect 256792 63504 256844 63510
rect 256698 63472 256754 63481
rect 204260 63436 204312 63442
rect 342260 63504 342312 63510
rect 256792 63446 256844 63452
rect 342258 63472 342260 63481
rect 342312 63472 342314 63481
rect 256698 63407 256700 63416
rect 204260 63378 204312 63384
rect 256752 63407 256754 63416
rect 256700 63378 256752 63384
rect 256804 62665 256832 63446
rect 342258 63407 342314 63416
rect 342352 63436 342404 63442
rect 342352 63378 342404 63384
rect 342364 62665 342392 63378
rect 256790 62656 256846 62665
rect 256790 62591 256846 62600
rect 342350 62656 342406 62665
rect 342350 62591 342406 62600
rect 256792 62076 256844 62082
rect 256792 62018 256844 62024
rect 342260 62076 342312 62082
rect 342260 62018 342312 62024
rect 198740 62008 198792 62014
rect 198740 61950 198792 61956
rect 256700 62008 256752 62014
rect 256700 61950 256752 61956
rect 256712 61849 256740 61950
rect 256698 61840 256754 61849
rect 256698 61775 256754 61784
rect 256804 61033 256832 62018
rect 342272 61849 342300 62018
rect 342352 62008 342404 62014
rect 342352 61950 342404 61956
rect 342258 61840 342314 61849
rect 342258 61775 342314 61784
rect 342364 61033 342392 61950
rect 256790 61024 256846 61033
rect 256790 60959 256846 60968
rect 342350 61024 342406 61033
rect 342350 60959 342406 60968
rect 256792 60716 256844 60722
rect 256792 60658 256844 60664
rect 342260 60716 342312 60722
rect 342260 60658 342312 60664
rect 191840 60648 191892 60654
rect 191840 60590 191892 60596
rect 256700 60648 256752 60654
rect 256700 60590 256752 60596
rect 256712 60353 256740 60590
rect 256698 60344 256754 60353
rect 256698 60279 256754 60288
rect 256804 59537 256832 60658
rect 342272 60353 342300 60658
rect 342352 60648 342404 60654
rect 342352 60590 342404 60596
rect 342258 60344 342314 60353
rect 342258 60279 342314 60288
rect 342364 59537 342392 60590
rect 256790 59528 256846 59537
rect 256790 59463 256846 59472
rect 342350 59528 342406 59537
rect 342350 59463 342406 59472
rect 186320 59356 186372 59362
rect 186320 59298 186372 59304
rect 256700 59356 256752 59362
rect 256700 59298 256752 59304
rect 342260 59356 342312 59362
rect 342260 59298 342312 59304
rect 256712 58721 256740 59298
rect 342272 58721 342300 59298
rect 256698 58712 256754 58721
rect 256698 58647 256754 58656
rect 342258 58712 342314 58721
rect 342258 58647 342314 58656
rect 256792 57928 256844 57934
rect 256698 57896 256754 57905
rect 183560 57860 183612 57866
rect 342260 57928 342312 57934
rect 256792 57870 256844 57876
rect 342258 57896 342260 57905
rect 342312 57896 342314 57905
rect 256698 57831 256700 57840
rect 183560 57802 183612 57808
rect 256752 57831 256754 57840
rect 256700 57802 256752 57808
rect 256804 57089 256832 57870
rect 342258 57831 342314 57840
rect 342352 57860 342404 57866
rect 342352 57802 342404 57808
rect 342364 57089 342392 57802
rect 256790 57080 256846 57089
rect 256790 57015 256846 57024
rect 342350 57080 342406 57089
rect 342350 57015 342406 57024
rect 256792 56568 256844 56574
rect 256792 56510 256844 56516
rect 342260 56568 342312 56574
rect 342260 56510 342312 56516
rect 176660 56500 176712 56506
rect 176660 56442 176712 56448
rect 256700 56500 256752 56506
rect 256700 56442 256752 56448
rect 256712 56273 256740 56442
rect 256698 56264 256754 56273
rect 256698 56199 256754 56208
rect 256804 55457 256832 56510
rect 342272 56273 342300 56510
rect 342352 56500 342404 56506
rect 342352 56442 342404 56448
rect 342258 56264 342314 56273
rect 342258 56199 342314 56208
rect 342364 55457 342392 56442
rect 256790 55448 256846 55457
rect 256790 55383 256846 55392
rect 342350 55448 342406 55457
rect 342350 55383 342406 55392
rect 171140 55208 171192 55214
rect 171140 55150 171192 55156
rect 256700 55208 256752 55214
rect 256700 55150 256752 55156
rect 342260 55208 342312 55214
rect 342260 55150 342312 55156
rect 256712 54641 256740 55150
rect 342272 54641 342300 55150
rect 256698 54632 256754 54641
rect 256698 54567 256754 54576
rect 342258 54632 342314 54641
rect 342258 54567 342314 54576
rect 256698 53816 256754 53825
rect 342258 53816 342314 53825
rect 256698 53751 256754 53760
rect 256792 53780 256844 53786
rect 256712 53718 256740 53751
rect 342258 53751 342260 53760
rect 256792 53722 256844 53728
rect 342312 53751 342314 53760
rect 342260 53722 342312 53728
rect 168380 53712 168432 53718
rect 168380 53654 168432 53660
rect 256700 53712 256752 53718
rect 256700 53654 256752 53660
rect 256804 53145 256832 53722
rect 342352 53712 342404 53718
rect 342352 53654 342404 53660
rect 342364 53145 342392 53654
rect 256790 53136 256846 53145
rect 256790 53071 256846 53080
rect 342350 53136 342406 53145
rect 342350 53071 342406 53080
rect 256792 52420 256844 52426
rect 256792 52362 256844 52368
rect 342260 52420 342312 52426
rect 342260 52362 342312 52368
rect 161480 52352 161532 52358
rect 256700 52352 256752 52358
rect 161480 52294 161532 52300
rect 256698 52320 256700 52329
rect 256752 52320 256754 52329
rect 256698 52255 256754 52264
rect 256804 51513 256832 52362
rect 342272 52329 342300 52362
rect 342352 52352 342404 52358
rect 342258 52320 342314 52329
rect 342352 52294 342404 52300
rect 342258 52255 342314 52264
rect 342364 51513 342392 52294
rect 256790 51504 256846 51513
rect 256790 51439 256846 51448
rect 342350 51504 342406 51513
rect 342350 51439 342406 51448
rect 256792 51060 256844 51066
rect 256792 51002 256844 51008
rect 342260 51060 342312 51066
rect 342260 51002 342312 51008
rect 155960 50992 156012 50998
rect 155960 50934 156012 50940
rect 256700 50992 256752 50998
rect 256700 50934 256752 50940
rect 256712 50697 256740 50934
rect 256698 50688 256754 50697
rect 256698 50623 256754 50632
rect 256804 49881 256832 51002
rect 342272 50697 342300 51002
rect 342352 50992 342404 50998
rect 342352 50934 342404 50940
rect 342258 50688 342314 50697
rect 342258 50623 342314 50632
rect 342364 49881 342392 50934
rect 256790 49872 256846 49881
rect 256790 49807 256846 49816
rect 342350 49872 342406 49881
rect 342350 49807 342406 49816
rect 149060 49700 149112 49706
rect 149060 49642 149112 49648
rect 256700 49700 256752 49706
rect 256700 49642 256752 49648
rect 342260 49700 342312 49706
rect 342260 49642 342312 49648
rect 256712 49065 256740 49642
rect 342272 49065 342300 49642
rect 256698 49056 256754 49065
rect 256698 48991 256754 49000
rect 342258 49056 342314 49065
rect 342258 48991 342314 49000
rect 256792 48272 256844 48278
rect 256698 48240 256754 48249
rect 146300 48204 146352 48210
rect 342260 48272 342312 48278
rect 256792 48214 256844 48220
rect 342258 48240 342260 48249
rect 342312 48240 342314 48249
rect 256698 48175 256700 48184
rect 146300 48146 146352 48152
rect 256752 48175 256754 48184
rect 256700 48146 256752 48152
rect 256804 47433 256832 48214
rect 342258 48175 342314 48184
rect 342352 48204 342404 48210
rect 342352 48146 342404 48152
rect 342364 47433 342392 48146
rect 256790 47424 256846 47433
rect 256790 47359 256846 47368
rect 342350 47424 342406 47433
rect 342350 47359 342406 47368
rect 256792 46912 256844 46918
rect 256792 46854 256844 46860
rect 342260 46912 342312 46918
rect 342260 46854 342312 46860
rect 140780 46844 140832 46850
rect 140780 46786 140832 46792
rect 256700 46844 256752 46850
rect 256700 46786 256752 46792
rect 256712 46753 256740 46786
rect 256698 46744 256754 46753
rect 256698 46679 256754 46688
rect 256804 45937 256832 46854
rect 342272 46753 342300 46854
rect 358096 46850 358124 438262
rect 359280 389836 359332 389842
rect 359280 389778 359332 389784
rect 358820 384600 358872 384606
rect 358820 384542 358872 384548
rect 358832 314265 358860 384542
rect 358912 384532 358964 384538
rect 358912 384474 358964 384480
rect 358924 315489 358952 384474
rect 359004 384464 359056 384470
rect 359004 384406 359056 384412
rect 359016 316985 359044 384406
rect 359096 384396 359148 384402
rect 359096 384338 359148 384344
rect 359108 318345 359136 384338
rect 359188 384328 359240 384334
rect 359188 384270 359240 384276
rect 359200 319977 359228 384270
rect 359292 379409 359320 389778
rect 359278 379400 359334 379409
rect 359278 379335 359334 379344
rect 359186 319968 359242 319977
rect 359186 319903 359242 319912
rect 359094 318336 359150 318345
rect 359094 318271 359150 318280
rect 359002 316976 359058 316985
rect 359002 316911 359058 316920
rect 358910 315480 358966 315489
rect 358910 315415 358966 315424
rect 358818 314256 358874 314265
rect 358818 314191 358874 314200
rect 379532 118590 379560 440014
rect 380912 385694 380940 440014
rect 381544 438524 381596 438530
rect 381544 438466 381596 438472
rect 380900 385688 380952 385694
rect 380900 385630 380952 385636
rect 379520 118584 379572 118590
rect 379520 118526 379572 118532
rect 342352 46844 342404 46850
rect 342352 46786 342404 46792
rect 358084 46844 358136 46850
rect 358084 46786 358136 46792
rect 342258 46744 342314 46753
rect 342258 46679 342314 46688
rect 342364 45937 342392 46786
rect 256790 45928 256846 45937
rect 256790 45863 256846 45872
rect 342350 45928 342406 45937
rect 342350 45863 342406 45872
rect 256792 45552 256844 45558
rect 256792 45494 256844 45500
rect 342352 45552 342404 45558
rect 342352 45494 342404 45500
rect 133880 45484 133932 45490
rect 133880 45426 133932 45432
rect 256700 45484 256752 45490
rect 256700 45426 256752 45432
rect 256712 45121 256740 45426
rect 256698 45112 256754 45121
rect 256698 45047 256754 45056
rect 256804 44305 256832 45494
rect 342260 45484 342312 45490
rect 342260 45426 342312 45432
rect 342272 45121 342300 45426
rect 342258 45112 342314 45121
rect 342258 45047 342314 45056
rect 342364 44305 342392 45494
rect 256790 44296 256846 44305
rect 256790 44231 256846 44240
rect 342350 44296 342406 44305
rect 342350 44231 342406 44240
rect 128360 44124 128412 44130
rect 128360 44066 128412 44072
rect 256700 44124 256752 44130
rect 256700 44066 256752 44072
rect 342260 44124 342312 44130
rect 342260 44066 342312 44072
rect 256712 43489 256740 44066
rect 342272 43489 342300 44066
rect 256698 43480 256754 43489
rect 256698 43415 256754 43424
rect 342258 43480 342314 43489
rect 342258 43415 342314 43424
rect 256792 42764 256844 42770
rect 256792 42706 256844 42712
rect 342260 42764 342312 42770
rect 342260 42706 342312 42712
rect 125600 42696 125652 42702
rect 256700 42696 256752 42702
rect 125600 42638 125652 42644
rect 256698 42664 256700 42673
rect 256752 42664 256754 42673
rect 256698 42599 256754 42608
rect 256804 41857 256832 42706
rect 342272 42673 342300 42706
rect 381556 42702 381584 438466
rect 382292 120086 382320 440014
rect 382924 438456 382976 438462
rect 382924 438398 382976 438404
rect 382280 120080 382332 120086
rect 382280 120022 382332 120028
rect 382936 42770 382964 438398
rect 383672 158778 383700 440014
rect 383660 158772 383712 158778
rect 383660 158714 383712 158720
rect 386432 118658 386460 440014
rect 386420 118652 386472 118658
rect 386420 118594 386472 118600
rect 387812 117230 387840 440014
rect 388444 438388 388496 438394
rect 388444 438330 388496 438336
rect 387800 117224 387852 117230
rect 387800 117166 387852 117172
rect 388456 45490 388484 438330
rect 388444 45484 388496 45490
rect 388444 45426 388496 45432
rect 382924 42764 382976 42770
rect 382924 42706 382976 42712
rect 342352 42696 342404 42702
rect 342258 42664 342314 42673
rect 342352 42638 342404 42644
rect 381544 42696 381596 42702
rect 381544 42638 381596 42644
rect 342258 42599 342314 42608
rect 342364 41857 342392 42638
rect 256790 41848 256846 41857
rect 256790 41783 256846 41792
rect 342350 41848 342406 41857
rect 342350 41783 342406 41792
rect 256792 41404 256844 41410
rect 256792 41346 256844 41352
rect 342260 41404 342312 41410
rect 342260 41346 342312 41352
rect 118700 41336 118752 41342
rect 118700 41278 118752 41284
rect 256700 41336 256752 41342
rect 256700 41278 256752 41284
rect 256712 41041 256740 41278
rect 256698 41032 256754 41041
rect 256698 40967 256754 40976
rect 256804 40361 256832 41346
rect 342272 41041 342300 41346
rect 389192 41342 389220 440014
rect 389824 437572 389876 437578
rect 389824 437514 389876 437520
rect 389836 41410 389864 437514
rect 390572 437510 390600 440014
rect 389916 437504 389968 437510
rect 389916 437446 389968 437452
rect 390560 437504 390612 437510
rect 390560 437446 390612 437452
rect 389928 92410 389956 437446
rect 389916 92404 389968 92410
rect 389916 92346 389968 92352
rect 391952 66162 391980 440014
rect 392584 438252 392636 438258
rect 392584 438194 392636 438200
rect 392596 106214 392624 438194
rect 393516 437578 393544 440014
rect 393964 438184 394016 438190
rect 393964 438126 394016 438132
rect 393504 437572 393556 437578
rect 393504 437514 393556 437520
rect 393976 107574 394004 438126
rect 393964 107568 394016 107574
rect 393964 107510 394016 107516
rect 392584 106208 392636 106214
rect 392584 106150 392636 106156
rect 394712 92478 394740 440014
rect 395344 438592 395396 438598
rect 395344 438534 395396 438540
rect 395356 95198 395384 438534
rect 395344 95192 395396 95198
rect 395344 95134 395396 95140
rect 394700 92472 394752 92478
rect 394700 92414 394752 92420
rect 396092 67522 396120 440014
rect 397932 438530 397960 440014
rect 397920 438524 397972 438530
rect 397920 438466 397972 438472
rect 398852 93770 398880 440014
rect 399484 437504 399536 437510
rect 399484 437446 399536 437452
rect 398840 93764 398892 93770
rect 398840 93706 398892 93712
rect 399496 69018 399524 437446
rect 399484 69012 399536 69018
rect 399484 68954 399536 68960
rect 400232 67590 400260 440014
rect 402348 438462 402376 440014
rect 402336 438456 402388 438462
rect 402336 438398 402388 438404
rect 402992 93838 403020 440014
rect 405292 437510 405320 440014
rect 405280 437504 405332 437510
rect 405280 437446 405332 437452
rect 402980 93832 403032 93838
rect 402980 93774 403032 93780
rect 400220 67584 400272 67590
rect 400220 67526 400272 67532
rect 396080 67516 396132 67522
rect 396080 67458 396132 67464
rect 391940 66156 391992 66162
rect 391940 66098 391992 66104
rect 405752 44130 405780 440014
rect 408512 438598 408540 440014
rect 408500 438592 408552 438598
rect 408500 438534 408552 438540
rect 409892 70310 409920 440014
rect 409880 70304 409932 70310
rect 409880 70246 409932 70252
rect 411272 45558 411300 440014
rect 412652 96558 412680 440014
rect 413284 438456 413336 438462
rect 413284 438398 413336 438404
rect 412640 96552 412692 96558
rect 412640 96494 412692 96500
rect 413296 71670 413324 438398
rect 413284 71664 413336 71670
rect 413284 71606 413336 71612
rect 414032 70378 414060 440014
rect 415596 438394 415624 440014
rect 415584 438388 415636 438394
rect 415584 438330 415636 438336
rect 416792 96626 416820 440014
rect 417424 438388 417476 438394
rect 417424 438330 417476 438336
rect 416780 96620 416832 96626
rect 416780 96562 416832 96568
rect 417436 73098 417464 438330
rect 417424 73092 417476 73098
rect 417424 73034 417476 73040
rect 418172 71738 418200 440014
rect 420012 438326 420040 440014
rect 420000 438320 420052 438326
rect 420000 438262 420052 438268
rect 420932 97918 420960 440014
rect 422956 438462 422984 440014
rect 422944 438456 422996 438462
rect 422944 438398 422996 438404
rect 420920 97912 420972 97918
rect 420920 97854 420972 97860
rect 418160 71732 418212 71738
rect 418160 71674 418212 71680
rect 414020 70372 414072 70378
rect 414020 70314 414072 70320
rect 423692 46918 423720 440014
rect 425072 97986 425100 440014
rect 427372 438394 427400 440014
rect 427360 438388 427412 438394
rect 427360 438330 427412 438336
rect 425060 97980 425112 97986
rect 425060 97922 425112 97928
rect 427832 48210 427860 440014
rect 430592 99346 430620 440014
rect 430580 99340 430632 99346
rect 430580 99282 430632 99288
rect 431972 73166 432000 440014
rect 431960 73160 432012 73166
rect 431960 73102 432012 73108
rect 433352 48278 433380 440014
rect 434732 100638 434760 440014
rect 434720 100632 434772 100638
rect 434720 100574 434772 100580
rect 436112 74526 436140 440014
rect 436100 74520 436152 74526
rect 436100 74462 436152 74468
rect 437492 49706 437520 440014
rect 438872 100706 438900 440014
rect 438860 100700 438912 100706
rect 438860 100642 438912 100648
rect 440252 75818 440280 440014
rect 440240 75812 440292 75818
rect 440240 75754 440292 75760
rect 441632 50998 441660 440014
rect 443012 102066 443040 440014
rect 445036 437510 445064 440014
rect 443644 437504 443696 437510
rect 443644 437446 443696 437452
rect 445024 437504 445076 437510
rect 445024 437446 445076 437452
rect 443000 102060 443052 102066
rect 443000 102002 443052 102008
rect 443656 75886 443684 437446
rect 443644 75880 443696 75886
rect 443644 75822 443696 75828
rect 445772 51066 445800 440014
rect 446404 438388 446456 438394
rect 446404 438330 446456 438336
rect 446416 60654 446444 438330
rect 447152 102134 447180 440014
rect 447140 102128 447192 102134
rect 447140 102070 447192 102076
rect 448532 77178 448560 440014
rect 448520 77172 448572 77178
rect 448520 77114 448572 77120
rect 446404 60648 446456 60654
rect 446404 60590 446456 60596
rect 449912 52358 449940 440014
rect 450544 438320 450596 438326
rect 450544 438262 450596 438268
rect 450556 60722 450584 438262
rect 452672 103426 452700 440014
rect 453304 438524 453356 438530
rect 453304 438466 453356 438472
rect 452660 103420 452712 103426
rect 452660 103362 452712 103368
rect 453316 79966 453344 438466
rect 453304 79960 453356 79966
rect 453304 79902 453356 79908
rect 454052 77246 454080 440014
rect 454040 77240 454092 77246
rect 454040 77182 454092 77188
rect 450544 60716 450596 60722
rect 450544 60658 450596 60664
rect 455432 52426 455460 440014
rect 456812 103494 456840 440014
rect 456800 103488 456852 103494
rect 456800 103430 456852 103436
rect 458192 78674 458220 440014
rect 458180 78668 458232 78674
rect 458180 78610 458232 78616
rect 459572 53718 459600 440014
rect 460204 438456 460256 438462
rect 460204 438398 460256 438404
rect 460216 62014 460244 438398
rect 460952 104854 460980 440014
rect 461584 438660 461636 438666
rect 461584 438602 461636 438608
rect 460940 104848 460992 104854
rect 460940 104790 460992 104796
rect 461596 82754 461624 438602
rect 462608 438530 462636 440014
rect 462596 438524 462648 438530
rect 462596 438466 462648 438472
rect 461584 82748 461636 82754
rect 461584 82690 461636 82696
rect 460204 62008 460256 62014
rect 460204 61950 460256 61956
rect 463712 53786 463740 440014
rect 464344 438524 464396 438530
rect 464344 438466 464396 438472
rect 464356 62082 464384 438466
rect 465092 106282 465120 440014
rect 465724 438728 465776 438734
rect 465724 438670 465776 438676
rect 465080 106276 465132 106282
rect 465080 106218 465132 106224
rect 465736 85474 465764 438670
rect 465724 85468 465776 85474
rect 465724 85410 465776 85416
rect 466472 80034 466500 440014
rect 466460 80028 466512 80034
rect 466460 79970 466512 79976
rect 464344 62076 464396 62082
rect 464344 62018 464396 62024
rect 467852 55214 467880 440014
rect 468484 438592 468536 438598
rect 468484 438534 468536 438540
rect 468496 63442 468524 438534
rect 469968 438258 469996 440014
rect 469956 438252 470008 438258
rect 469956 438194 470008 438200
rect 470612 81326 470640 440014
rect 470600 81320 470652 81326
rect 470600 81262 470652 81268
rect 468484 63436 468536 63442
rect 468484 63378 468536 63384
rect 471992 56506 472020 440014
rect 472624 438252 472676 438258
rect 472624 438194 472676 438200
rect 472636 63510 472664 438194
rect 474384 438190 474412 440014
rect 474372 438184 474424 438190
rect 474372 438126 474424 438132
rect 475384 438184 475436 438190
rect 475384 438126 475436 438132
rect 475396 64870 475424 438126
rect 476132 81394 476160 440014
rect 476120 81388 476172 81394
rect 476120 81330 476172 81336
rect 475384 64864 475436 64870
rect 475384 64806 475436 64812
rect 472624 63504 472676 63510
rect 472624 63446 472676 63452
rect 477512 56574 477540 440014
rect 478892 107642 478920 440014
rect 480364 438666 480392 440014
rect 480352 438660 480404 438666
rect 480352 438602 480404 438608
rect 478880 107636 478932 107642
rect 478880 107578 478932 107584
rect 481652 57866 481680 440014
rect 482284 438660 482336 438666
rect 482284 438602 482336 438608
rect 482296 66230 482324 438602
rect 483032 108934 483060 440014
rect 483020 108928 483072 108934
rect 483020 108870 483072 108876
rect 484412 82822 484440 440014
rect 484400 82816 484452 82822
rect 484400 82758 484452 82764
rect 482284 66224 482336 66230
rect 482284 66166 482336 66172
rect 485792 57934 485820 440014
rect 487632 437510 487660 440014
rect 486424 437504 486476 437510
rect 486424 437446 486476 437452
rect 487620 437504 487672 437510
rect 487620 437446 487672 437452
rect 486436 109002 486464 437446
rect 486424 108996 486476 109002
rect 486424 108938 486476 108944
rect 488552 84182 488580 440014
rect 488540 84176 488592 84182
rect 488540 84118 488592 84124
rect 489932 59362 489960 440014
rect 492048 437510 492076 440014
rect 490564 437504 490616 437510
rect 490564 437446 490616 437452
rect 492036 437504 492088 437510
rect 492036 437446 492088 437452
rect 490576 110430 490604 437446
rect 490564 110424 490616 110430
rect 490564 110366 490616 110372
rect 492692 85542 492720 440014
rect 494992 438394 495020 440014
rect 494980 438388 495032 438394
rect 494980 438330 495032 438336
rect 496464 437510 496492 440014
rect 498212 438734 498240 440014
rect 498200 438728 498252 438734
rect 498200 438670 498252 438676
rect 499592 438326 499620 440014
rect 499580 438320 499632 438326
rect 499580 438262 499632 438268
rect 500972 437578 501000 440014
rect 501604 438320 501656 438326
rect 501604 438262 501656 438268
rect 497464 437572 497516 437578
rect 497464 437514 497516 437520
rect 500960 437572 501012 437578
rect 500960 437514 501012 437520
rect 494704 437504 494756 437510
rect 494704 437446 494756 437452
rect 496452 437504 496504 437510
rect 496452 437446 496504 437452
rect 494716 111722 494744 437446
rect 497476 111790 497504 437514
rect 500224 437504 500276 437510
rect 500224 437446 500276 437452
rect 500236 113082 500264 437446
rect 501616 113150 501644 438262
rect 501604 113144 501656 113150
rect 501604 113086 501656 113092
rect 500224 113076 500276 113082
rect 500224 113018 500276 113024
rect 497464 111784 497516 111790
rect 497464 111726 497516 111732
rect 494704 111716 494756 111722
rect 494704 111658 494756 111664
rect 502352 86902 502380 440014
rect 503824 438462 503852 440014
rect 503812 438456 503864 438462
rect 503812 438398 503864 438404
rect 504364 438456 504416 438462
rect 504364 438398 504416 438404
rect 504376 114510 504404 438398
rect 505296 437510 505324 440014
rect 505284 437504 505336 437510
rect 505284 437446 505336 437452
rect 504364 114504 504416 114510
rect 504364 114446 504416 114452
rect 506492 86970 506520 440014
rect 508240 438530 508268 440014
rect 508228 438524 508280 438530
rect 508228 438466 508280 438472
rect 508504 438388 508556 438394
rect 508504 438330 508556 438336
rect 508516 115870 508544 438330
rect 509712 438326 509740 440014
rect 509700 438320 509752 438326
rect 509700 438262 509752 438268
rect 508504 115864 508556 115870
rect 508504 115806 508556 115812
rect 510632 88262 510660 440014
rect 512656 438598 512684 440014
rect 512644 438592 512696 438598
rect 512644 438534 512696 438540
rect 514128 438462 514156 440014
rect 514116 438456 514168 438462
rect 514116 438398 514168 438404
rect 512644 438320 512696 438326
rect 512644 438262 512696 438268
rect 512656 115938 512684 438262
rect 512644 115932 512696 115938
rect 512644 115874 512696 115880
rect 514772 88330 514800 440014
rect 517072 438258 517100 440014
rect 518544 438394 518572 440014
rect 518532 438388 518584 438394
rect 518532 438330 518584 438336
rect 517060 438252 517112 438258
rect 517060 438194 517112 438200
rect 518164 438252 518216 438258
rect 518164 438194 518216 438200
rect 518176 117298 518204 438194
rect 520292 437510 520320 440014
rect 521672 438190 521700 440014
rect 523052 438326 523080 440014
rect 523040 438320 523092 438326
rect 523040 438262 523092 438268
rect 521660 438184 521712 438190
rect 521660 438126 521712 438132
rect 524432 437578 524460 440014
rect 525904 438666 525932 440014
rect 525892 438660 525944 438666
rect 525892 438602 525944 438608
rect 527376 438258 527404 440014
rect 527364 438252 527416 438258
rect 527364 438194 527416 438200
rect 520924 437572 520976 437578
rect 520924 437514 520976 437520
rect 524420 437572 524472 437578
rect 524420 437514 524472 437520
rect 519544 437504 519596 437510
rect 519544 437446 519596 437452
rect 520280 437504 520332 437510
rect 520280 437446 520332 437452
rect 518164 117292 518216 117298
rect 518164 117234 518216 117240
rect 519556 89690 519584 437446
rect 520936 90982 520964 437514
rect 528848 437510 528876 440014
rect 522304 437504 522356 437510
rect 522304 437446 522356 437452
rect 528836 437504 528888 437510
rect 528836 437446 528888 437452
rect 522316 91050 522344 437446
rect 548536 379506 548564 552298
rect 551296 431934 551324 552366
rect 555424 552288 555476 552294
rect 555424 552230 555476 552236
rect 554044 552220 554096 552226
rect 554044 552162 554096 552168
rect 554056 471986 554084 552162
rect 555436 525774 555464 552230
rect 556804 552152 556856 552158
rect 556804 552094 556856 552100
rect 555424 525768 555476 525774
rect 555424 525710 555476 525716
rect 554044 471980 554096 471986
rect 554044 471922 554096 471928
rect 551284 431928 551336 431934
rect 551284 431870 551336 431876
rect 548524 379500 548576 379506
rect 548524 379442 548576 379448
rect 556816 365702 556844 552094
rect 558184 552084 558236 552090
rect 558184 552026 558236 552032
rect 558196 419490 558224 552026
rect 580264 549296 580316 549302
rect 580264 549238 580316 549244
rect 579896 538212 579948 538218
rect 579896 538154 579948 538160
rect 579908 537849 579936 538154
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580276 484673 580304 549238
rect 580262 484664 580318 484673
rect 580262 484599 580318 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 431633 579844 431870
rect 579802 431624 579858 431633
rect 579802 431559 579858 431568
rect 558184 419484 558236 419490
rect 558184 419426 558236 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 556804 365696 556856 365702
rect 556804 365638 556856 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 522304 91044 522356 91050
rect 522304 90986 522356 90992
rect 520924 90976 520976 90982
rect 520924 90918 520976 90924
rect 519544 89684 519596 89690
rect 519544 89626 519596 89632
rect 514760 88324 514812 88330
rect 514760 88266 514812 88272
rect 510620 88256 510672 88262
rect 510620 88198 510672 88204
rect 506480 86964 506532 86970
rect 506480 86906 506532 86912
rect 502340 86896 502392 86902
rect 502340 86838 502392 86844
rect 492680 85536 492732 85542
rect 492680 85478 492732 85484
rect 489920 59356 489972 59362
rect 489920 59298 489972 59304
rect 485780 57928 485832 57934
rect 485780 57870 485832 57876
rect 481640 57860 481692 57866
rect 481640 57802 481692 57808
rect 477500 56568 477552 56574
rect 477500 56510 477552 56516
rect 471980 56500 472032 56506
rect 471980 56442 472032 56448
rect 467840 55208 467892 55214
rect 467840 55150 467892 55156
rect 463700 53780 463752 53786
rect 463700 53722 463752 53728
rect 459560 53712 459612 53718
rect 459560 53654 459612 53660
rect 455420 52420 455472 52426
rect 455420 52362 455472 52368
rect 449900 52352 449952 52358
rect 449900 52294 449952 52300
rect 445760 51060 445812 51066
rect 445760 51002 445812 51008
rect 441620 50992 441672 50998
rect 441620 50934 441672 50940
rect 437480 49700 437532 49706
rect 437480 49642 437532 49648
rect 433340 48272 433392 48278
rect 433340 48214 433392 48220
rect 427820 48204 427872 48210
rect 427820 48146 427872 48152
rect 423680 46912 423732 46918
rect 423680 46854 423732 46860
rect 411260 45552 411312 45558
rect 411260 45494 411312 45500
rect 405740 44124 405792 44130
rect 405740 44066 405792 44072
rect 389824 41404 389876 41410
rect 389824 41346 389876 41352
rect 342352 41336 342404 41342
rect 342352 41278 342404 41284
rect 389180 41336 389232 41342
rect 389180 41278 389232 41284
rect 342258 41032 342314 41041
rect 342258 40967 342314 40976
rect 342364 40361 342392 41278
rect 256790 40352 256846 40361
rect 256790 40287 256846 40296
rect 342350 40352 342406 40361
rect 342350 40287 342406 40296
rect 259472 40038 260406 40066
rect 260852 40038 261142 40066
rect 261220 40038 261970 40066
rect 262232 40038 262798 40066
rect 263152 40038 263534 40066
rect 263612 40038 264362 40066
rect 265084 40038 265190 40066
rect 265544 40038 265926 40066
rect 266464 40038 266754 40066
rect 267200 40038 267582 40066
rect 267752 40038 268410 40066
rect 124220 38412 124272 38418
rect 124220 38354 124272 38360
rect 120080 21684 120132 21690
rect 120080 21626 120132 21632
rect 113272 21616 113324 21622
rect 113272 21558 113324 21564
rect 113284 16574 113312 21558
rect 120092 16574 120120 21626
rect 124232 16574 124260 38354
rect 113284 16546 114048 16574
rect 120092 16546 120672 16574
rect 124232 16546 124720 16574
rect 113180 9240 113232 9246
rect 113180 9182 113232 9188
rect 112812 8152 112864 8158
rect 112812 8094 112864 8100
rect 112824 480 112852 8094
rect 114020 480 114048 16546
rect 118792 13456 118844 13462
rect 118792 13398 118844 13404
rect 114744 12164 114796 12170
rect 114744 12106 114796 12112
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 12106
rect 116400 8220 116452 8226
rect 116400 8162 116452 8168
rect 116412 480 116440 8162
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 117608 480 117636 3674
rect 118804 480 118832 13398
rect 119896 9240 119948 9246
rect 119896 9182 119948 9188
rect 119908 480 119936 9182
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 123024 16312 123076 16318
rect 123024 16254 123076 16260
rect 122288 13524 122340 13530
rect 122288 13466 122340 13472
rect 122300 480 122328 13466
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16254
rect 124692 480 124720 16546
rect 259472 9042 259500 40038
rect 260852 10334 260880 40038
rect 261220 26234 261248 40038
rect 260944 26206 261248 26234
rect 260944 11762 260972 26206
rect 262232 11830 262260 40038
rect 263152 26234 263180 40038
rect 262324 26206 263180 26234
rect 262324 13190 262352 26206
rect 262312 13184 262364 13190
rect 262312 13126 262364 13132
rect 262220 11824 262272 11830
rect 262220 11766 262272 11772
rect 260932 11756 260984 11762
rect 260932 11698 260984 11704
rect 260840 10328 260892 10334
rect 260840 10270 260892 10276
rect 259460 9036 259512 9042
rect 259460 8978 259512 8984
rect 263612 6526 263640 40038
rect 264980 37868 265032 37874
rect 264980 37810 265032 37816
rect 264992 13394 265020 37810
rect 264980 13388 265032 13394
rect 264980 13330 265032 13336
rect 265084 13326 265112 40038
rect 265544 37874 265572 40038
rect 265532 37868 265584 37874
rect 265532 37810 265584 37816
rect 266360 37868 266412 37874
rect 266360 37810 266412 37816
rect 265072 13320 265124 13326
rect 265072 13262 265124 13268
rect 266372 6662 266400 37810
rect 266360 6656 266412 6662
rect 266360 6598 266412 6604
rect 266464 6594 266492 40038
rect 267200 37874 267228 40038
rect 267188 37868 267240 37874
rect 267188 37810 267240 37816
rect 267752 9110 267780 40038
rect 269132 9178 269160 40052
rect 269224 40038 269974 40066
rect 270604 40038 270802 40066
rect 271248 40038 271538 40066
rect 271984 40038 272366 40066
rect 272904 40038 273194 40066
rect 273272 40038 273930 40066
rect 269224 10402 269252 40038
rect 270500 37868 270552 37874
rect 270500 37810 270552 37816
rect 270512 10538 270540 37810
rect 270500 10532 270552 10538
rect 270500 10474 270552 10480
rect 270604 10470 270632 40038
rect 271248 37874 271276 40038
rect 271236 37868 271288 37874
rect 271236 37810 271288 37816
rect 271880 36440 271932 36446
rect 271880 36382 271932 36388
rect 271892 10674 271920 36382
rect 271880 10668 271932 10674
rect 271880 10610 271932 10616
rect 271984 10606 272012 40038
rect 272904 36446 272932 40038
rect 272892 36440 272944 36446
rect 272892 36382 272944 36388
rect 271972 10600 272024 10606
rect 271972 10542 272024 10548
rect 270592 10464 270644 10470
rect 270592 10406 270644 10412
rect 269212 10396 269264 10402
rect 269212 10338 269264 10344
rect 269120 9172 269172 9178
rect 269120 9114 269172 9120
rect 267740 9104 267792 9110
rect 267740 9046 267792 9052
rect 266452 6588 266504 6594
rect 266452 6530 266504 6536
rect 263600 6520 263652 6526
rect 263600 6462 263652 6468
rect 273272 4826 273300 40038
rect 274640 37868 274692 37874
rect 274640 37810 274692 37816
rect 274652 4962 274680 37810
rect 274640 4956 274692 4962
rect 274640 4898 274692 4904
rect 274744 4894 274772 40052
rect 275296 40038 275586 40066
rect 276124 40038 276414 40066
rect 276768 40038 277150 40066
rect 277412 40038 277978 40066
rect 275296 37874 275324 40038
rect 275284 37868 275336 37874
rect 275284 37810 275336 37816
rect 276020 37868 276072 37874
rect 276020 37810 276072 37816
rect 276032 5098 276060 37810
rect 276020 5092 276072 5098
rect 276020 5034 276072 5040
rect 276124 5030 276152 40038
rect 276768 37874 276796 40038
rect 276756 37868 276808 37874
rect 276756 37810 276808 37816
rect 277412 5166 277440 40038
rect 278792 11898 278820 40052
rect 278884 40038 279542 40066
rect 280172 40038 280370 40066
rect 280448 40038 281198 40066
rect 281552 40038 281934 40066
rect 282104 40038 282762 40066
rect 282932 40038 283590 40066
rect 284312 40038 284418 40066
rect 284680 40038 285154 40066
rect 285692 40038 285982 40066
rect 286060 40038 286810 40066
rect 287072 40038 287546 40066
rect 287624 40038 288374 40066
rect 288452 40038 289202 40066
rect 289832 40038 289938 40066
rect 290016 40038 290766 40066
rect 291212 40038 291594 40066
rect 291856 40038 292422 40066
rect 292592 40038 293158 40066
rect 278884 11966 278912 40038
rect 278872 11960 278924 11966
rect 278872 11902 278924 11908
rect 278780 11892 278832 11898
rect 278780 11834 278832 11840
rect 280172 5234 280200 40038
rect 280448 26234 280476 40038
rect 280264 26206 280476 26234
rect 280264 12034 280292 26206
rect 280252 12028 280304 12034
rect 280252 11970 280304 11976
rect 281552 9314 281580 40038
rect 282104 26234 282132 40038
rect 281644 26206 282132 26234
rect 281644 12102 281672 26206
rect 282932 12170 282960 40038
rect 284312 13462 284340 40038
rect 284680 26234 284708 40038
rect 284404 26206 284708 26234
rect 284404 13530 284432 26206
rect 284392 13524 284444 13530
rect 284392 13466 284444 13472
rect 284300 13456 284352 13462
rect 284300 13398 284352 13404
rect 282920 12164 282972 12170
rect 282920 12106 282972 12112
rect 281632 12096 281684 12102
rect 281632 12038 281684 12044
rect 281540 9308 281592 9314
rect 281540 9250 281592 9256
rect 285692 6254 285720 40038
rect 286060 26234 286088 40038
rect 285784 26206 286088 26234
rect 285784 13122 285812 26206
rect 285772 13116 285824 13122
rect 285772 13058 285824 13064
rect 287072 7614 287100 40038
rect 287624 26234 287652 40038
rect 287164 26206 287652 26234
rect 287164 15910 287192 26206
rect 288452 15978 288480 40038
rect 289832 16046 289860 40038
rect 290016 26234 290044 40038
rect 289924 26206 290044 26234
rect 289924 16114 289952 26206
rect 291212 16182 291240 40038
rect 291856 26234 291884 40038
rect 291304 26206 291884 26234
rect 291304 17542 291332 26206
rect 292592 17610 292620 40038
rect 292580 17604 292632 17610
rect 292580 17546 292632 17552
rect 291292 17536 291344 17542
rect 291292 17478 291344 17484
rect 291200 16176 291252 16182
rect 291200 16118 291252 16124
rect 289912 16108 289964 16114
rect 289912 16050 289964 16056
rect 289820 16040 289872 16046
rect 289820 15982 289872 15988
rect 288440 15972 288492 15978
rect 288440 15914 288492 15920
rect 287152 15904 287204 15910
rect 287152 15846 287204 15852
rect 287060 7608 287112 7614
rect 287060 7550 287112 7556
rect 293972 6322 294000 40052
rect 294064 40038 294814 40066
rect 295352 40038 295550 40066
rect 295904 40038 296378 40066
rect 296732 40038 297206 40066
rect 297468 40038 297942 40066
rect 298112 40038 298770 40066
rect 299492 40038 299598 40066
rect 299952 40038 300426 40066
rect 300872 40038 301162 40066
rect 301516 40038 301990 40066
rect 302252 40038 302818 40066
rect 302988 40038 303554 40066
rect 303632 40038 304382 40066
rect 305012 40038 305210 40066
rect 305472 40038 305946 40066
rect 306392 40038 306774 40066
rect 307312 40038 307602 40066
rect 307772 40038 308430 40066
rect 294064 6390 294092 40038
rect 295352 6458 295380 40038
rect 295904 26234 295932 40038
rect 295444 26206 295932 26234
rect 295444 13258 295472 26206
rect 296732 14482 296760 40038
rect 297468 26234 297496 40038
rect 296824 26206 297496 26234
rect 296824 14550 296852 26206
rect 298112 14618 298140 40038
rect 299492 14686 299520 40038
rect 299952 26234 299980 40038
rect 299584 26206 299980 26234
rect 299584 14754 299612 26206
rect 300872 14822 300900 40038
rect 301516 26234 301544 40038
rect 300964 26206 301544 26234
rect 300964 16250 300992 26206
rect 300952 16244 301004 16250
rect 300952 16186 301004 16192
rect 300860 14816 300912 14822
rect 300860 14758 300912 14764
rect 299572 14748 299624 14754
rect 299572 14690 299624 14696
rect 299480 14680 299532 14686
rect 299480 14622 299532 14628
rect 298100 14612 298152 14618
rect 298100 14554 298152 14560
rect 296812 14544 296864 14550
rect 296812 14486 296864 14492
rect 296720 14476 296772 14482
rect 296720 14418 296772 14424
rect 295432 13252 295484 13258
rect 295432 13194 295484 13200
rect 302252 7682 302280 40038
rect 302988 26234 303016 40038
rect 302344 26206 303016 26234
rect 302344 7750 302372 26206
rect 303632 7818 303660 40038
rect 305012 7886 305040 40038
rect 305472 26234 305500 40038
rect 305104 26206 305500 26234
rect 305104 7954 305132 26206
rect 306392 8022 306420 40038
rect 307312 26234 307340 40038
rect 306484 26206 307340 26234
rect 306484 8090 306512 26206
rect 307772 8158 307800 40038
rect 309152 8226 309180 40052
rect 309244 40038 309994 40066
rect 310532 40038 310822 40066
rect 311176 40038 311558 40066
rect 312004 40038 312386 40066
rect 309244 9246 309272 40038
rect 310532 16318 310560 40038
rect 311176 26234 311204 40038
rect 310624 26206 311204 26234
rect 310624 17270 310652 26206
rect 312004 19990 312032 40038
rect 313200 38010 313228 40052
rect 313292 40038 313950 40066
rect 313188 38004 313240 38010
rect 313188 37946 313240 37952
rect 311992 19984 312044 19990
rect 311992 19926 312044 19932
rect 310612 17264 310664 17270
rect 310612 17206 310664 17212
rect 310520 16312 310572 16318
rect 310520 16254 310572 16260
rect 309232 9240 309284 9246
rect 309232 9182 309284 9188
rect 309140 8220 309192 8226
rect 309140 8162 309192 8168
rect 307760 8152 307812 8158
rect 307760 8094 307812 8100
rect 306472 8084 306524 8090
rect 306472 8026 306524 8032
rect 306380 8016 306432 8022
rect 306380 7958 306432 7964
rect 305092 7948 305144 7954
rect 305092 7890 305144 7896
rect 305000 7880 305052 7886
rect 305000 7822 305052 7828
rect 303620 7812 303672 7818
rect 303620 7754 303672 7760
rect 302332 7744 302384 7750
rect 302332 7686 302384 7692
rect 302240 7676 302292 7682
rect 302240 7618 302292 7624
rect 295340 6452 295392 6458
rect 295340 6394 295392 6400
rect 294052 6384 294104 6390
rect 294052 6326 294104 6332
rect 293960 6316 294012 6322
rect 293960 6258 294012 6264
rect 285680 6248 285732 6254
rect 285680 6190 285732 6196
rect 280160 5228 280212 5234
rect 280160 5170 280212 5176
rect 277400 5160 277452 5166
rect 277400 5102 277452 5108
rect 276112 5024 276164 5030
rect 276112 4966 276164 4972
rect 274732 4888 274784 4894
rect 274732 4830 274784 4836
rect 273260 4820 273312 4826
rect 273260 4762 273312 4768
rect 313292 3534 313320 40038
rect 314764 38078 314792 40052
rect 315132 40038 315606 40066
rect 314752 38072 314804 38078
rect 314752 38014 314804 38020
rect 315132 26234 315160 40038
rect 316420 38214 316448 40052
rect 316512 40038 317170 40066
rect 316408 38208 316460 38214
rect 316408 38150 316460 38156
rect 316512 26234 316540 40038
rect 317984 38146 318012 40052
rect 318834 40038 318932 40066
rect 317972 38140 318024 38146
rect 317972 38082 318024 38088
rect 318800 38004 318852 38010
rect 318800 37946 318852 37952
rect 314764 26206 315160 26234
rect 316144 26206 316540 26234
rect 314764 3602 314792 26206
rect 316144 3670 316172 26206
rect 318812 17338 318840 37946
rect 318904 21418 318932 40038
rect 319272 40038 319562 40066
rect 320284 40038 320390 40066
rect 320928 40038 321218 40066
rect 321664 40038 321954 40066
rect 322400 40038 322782 40066
rect 322952 40038 323610 40066
rect 324332 40038 324438 40066
rect 324608 40038 325174 40066
rect 325712 40038 326002 40066
rect 326080 40038 326830 40066
rect 327092 40038 327566 40066
rect 327644 40038 328394 40066
rect 328472 40038 329222 40066
rect 319272 38010 319300 40038
rect 319260 38004 319312 38010
rect 319260 37946 319312 37952
rect 320180 38004 320232 38010
rect 320180 37946 320232 37952
rect 318892 21412 318944 21418
rect 318892 21354 318944 21360
rect 320192 17474 320220 37946
rect 320180 17468 320232 17474
rect 320180 17410 320232 17416
rect 320284 17406 320312 40038
rect 320824 38072 320876 38078
rect 320824 38014 320876 38020
rect 320272 17400 320324 17406
rect 320272 17342 320324 17348
rect 318800 17332 318852 17338
rect 318800 17274 318852 17280
rect 320836 3738 320864 38014
rect 320928 38010 320956 40038
rect 320916 38004 320968 38010
rect 320916 37946 320968 37952
rect 321560 35896 321612 35902
rect 321560 35838 321612 35844
rect 321572 18698 321600 35838
rect 321560 18692 321612 18698
rect 321560 18634 321612 18640
rect 321664 18630 321692 40038
rect 322204 38072 322256 38078
rect 322204 38014 322256 38020
rect 321652 18624 321704 18630
rect 321652 18566 321704 18572
rect 320824 3732 320876 3738
rect 320824 3674 320876 3680
rect 316132 3664 316184 3670
rect 316132 3606 316184 3612
rect 314752 3596 314804 3602
rect 314752 3538 314804 3544
rect 313280 3528 313332 3534
rect 313280 3470 313332 3476
rect 322216 3466 322244 38014
rect 322400 35902 322428 40038
rect 322388 35896 322440 35902
rect 322388 35838 322440 35844
rect 322952 18766 322980 40038
rect 324332 18834 324360 40038
rect 324608 26234 324636 40038
rect 324424 26206 324636 26234
rect 324424 18902 324452 26206
rect 325712 18970 325740 40038
rect 326080 26234 326108 40038
rect 325804 26206 326108 26234
rect 325804 20058 325832 26206
rect 327092 20126 327120 40038
rect 327644 26234 327672 40038
rect 327184 26206 327672 26234
rect 327184 20194 327212 26206
rect 328472 20262 328500 40038
rect 329944 20330 329972 40052
rect 330772 38282 330800 40052
rect 331324 40038 331614 40066
rect 330760 38276 330812 38282
rect 330760 38218 330812 38224
rect 331324 21486 331352 40038
rect 332428 38350 332456 40052
rect 332612 40038 333178 40066
rect 334014 40038 334112 40066
rect 332416 38344 332468 38350
rect 332416 38286 332468 38292
rect 332612 21554 332640 40038
rect 334084 21622 334112 40038
rect 334820 38010 334848 40052
rect 335464 40038 335570 40066
rect 334808 38004 334860 38010
rect 334808 37946 334860 37952
rect 335464 21690 335492 40038
rect 336384 38418 336412 40052
rect 336372 38412 336424 38418
rect 336372 38354 336424 38360
rect 337212 38078 337240 40052
rect 337200 38072 337252 38078
rect 337200 38014 337252 38020
rect 337948 37942 337976 40052
rect 338132 40038 338790 40066
rect 339512 40038 339618 40066
rect 337936 37936 337988 37942
rect 337936 37878 337988 37884
rect 335452 21684 335504 21690
rect 335452 21626 335504 21632
rect 334072 21616 334124 21622
rect 334072 21558 334124 21564
rect 332600 21548 332652 21554
rect 332600 21490 332652 21496
rect 331312 21480 331364 21486
rect 331312 21422 331364 21428
rect 329932 20324 329984 20330
rect 329932 20266 329984 20272
rect 328460 20256 328512 20262
rect 328460 20198 328512 20204
rect 327172 20188 327224 20194
rect 327172 20130 327224 20136
rect 327080 20120 327132 20126
rect 327080 20062 327132 20068
rect 325792 20052 325844 20058
rect 325792 19994 325844 20000
rect 325700 18964 325752 18970
rect 325700 18906 325752 18912
rect 324412 18896 324464 18902
rect 324412 18838 324464 18844
rect 324320 18828 324372 18834
rect 324320 18770 324372 18776
rect 322940 18760 322992 18766
rect 322940 18702 322992 18708
rect 338132 8974 338160 40038
rect 338120 8968 338172 8974
rect 338120 8910 338172 8916
rect 339512 6186 339540 40038
rect 339500 6180 339552 6186
rect 339500 6122 339552 6128
rect 322204 3460 322256 3466
rect 322204 3402 322256 3408
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 376942 548664 376998 548720
rect 251822 499024 251878 499080
rect 251914 495216 251970 495272
rect 251270 486920 251326 486976
rect 251362 485596 251364 485616
rect 251364 485596 251416 485616
rect 251416 485596 251418 485616
rect 251362 485560 251418 485596
rect 251730 485016 251786 485072
rect 251730 483928 251786 483984
rect 251730 481208 251786 481264
rect 252006 491136 252062 491192
rect 251914 490592 251970 490648
rect 251822 479440 251878 479496
rect 252466 499296 252522 499352
rect 252466 497800 252522 497856
rect 252466 496748 252468 496768
rect 252468 496748 252520 496768
rect 252520 496748 252522 496768
rect 252466 496712 252522 496748
rect 252374 496168 252430 496224
rect 252466 493992 252522 494048
rect 252374 493448 252430 493504
rect 252466 492088 252522 492144
rect 252466 489504 252522 489560
rect 252466 488452 252468 488472
rect 252468 488452 252520 488472
rect 252520 488452 252522 488472
rect 252466 488416 252522 488452
rect 252098 487872 252154 487928
rect 376942 546080 376998 546136
rect 376850 543496 376906 543552
rect 377402 540912 377458 540968
rect 376942 538328 376998 538384
rect 376942 535880 376998 535936
rect 376942 533296 376998 533352
rect 376942 528128 376998 528184
rect 376942 525544 376998 525600
rect 376942 523096 376998 523152
rect 376942 517928 376998 517984
rect 376942 515344 376998 515400
rect 376942 512760 376998 512816
rect 376942 510176 376998 510232
rect 377494 530712 377550 530768
rect 377402 494944 377458 495000
rect 376942 492360 376998 492416
rect 376942 489776 376998 489832
rect 376942 487212 376998 487248
rect 376942 487192 376944 487212
rect 376944 487192 376996 487212
rect 376996 487192 376998 487212
rect 252466 482840 252522 482896
rect 252374 482296 252430 482352
rect 377218 482160 377274 482216
rect 252466 479984 252522 480040
rect 377034 479576 377090 479632
rect 252006 478488 252062 478544
rect 251914 477400 251970 477456
rect 376942 476992 376998 477048
rect 251730 476720 251786 476776
rect 252466 475632 252522 475688
rect 377586 520512 377642 520568
rect 377678 507728 377734 507784
rect 377770 505144 377826 505200
rect 377862 502560 377918 502616
rect 377494 484608 377550 484664
rect 377954 499976 378010 500032
rect 378046 497392 378102 497448
rect 252466 474408 252522 474464
rect 376942 474408 376998 474464
rect 251914 473864 251970 473920
rect 251546 472912 251602 472968
rect 376942 471824 376998 471880
rect 252466 471416 252522 471472
rect 252466 470736 252522 470792
rect 252466 469240 252522 469296
rect 376942 469240 376998 469296
rect 252374 468152 252430 468208
rect 251546 467200 251602 467256
rect 251270 464480 251326 464536
rect 252282 465432 252338 465488
rect 252190 463664 252246 463720
rect 252006 462576 252062 462632
rect 251914 461080 251970 461136
rect 68742 386280 68798 386336
rect 71318 386280 71374 386336
rect 78494 386316 78496 386336
rect 78496 386316 78548 386336
rect 78548 386316 78550 386336
rect 78494 386280 78550 386316
rect 89166 386316 89168 386336
rect 89168 386316 89220 386336
rect 89220 386316 89222 386336
rect 89166 386280 89222 386316
rect 93766 386280 93822 386336
rect 96526 386280 96582 386336
rect 99286 386280 99342 386336
rect 102046 386280 102102 386336
rect 73894 385056 73950 385112
rect 77206 385056 77262 385112
rect 81070 385056 81126 385112
rect 83646 385092 83648 385112
rect 83648 385092 83700 385112
rect 83700 385092 83702 385112
rect 83646 385056 83702 385092
rect 106186 386280 106242 386336
rect 108946 386280 109002 386336
rect 111706 386280 111762 386336
rect 104806 385192 104862 385248
rect 117226 386280 117282 386336
rect 118606 386280 118662 386336
rect 124126 386280 124182 386336
rect 126886 386280 126942 386336
rect 133694 386316 133696 386336
rect 133696 386316 133748 386336
rect 133748 386316 133750 386336
rect 133694 386280 133750 386316
rect 86498 385056 86554 385112
rect 92110 385056 92166 385112
rect 114466 385056 114522 385112
rect 121366 385056 121422 385112
rect 128634 385056 128690 385112
rect 131026 385056 131082 385112
rect 136086 385056 136142 385112
rect 138478 386316 138480 386336
rect 138480 386316 138532 386336
rect 138532 386316 138534 386336
rect 138478 386280 138534 386316
rect 142066 386280 142122 386336
rect 143446 386280 143502 386336
rect 158534 386280 158590 386336
rect 159822 386280 159878 386336
rect 146206 385056 146262 385112
rect 170862 384104 170918 384160
rect 38290 336776 38346 336832
rect 38750 335552 38806 335608
rect 38382 333104 38438 333160
rect 38566 332560 38622 332616
rect 38474 309304 38530 309360
rect 38382 229744 38438 229800
rect 38658 327528 38714 327584
rect 39026 330384 39082 330440
rect 38842 329840 38898 329896
rect 38934 307808 38990 307864
rect 39118 308352 39174 308408
rect 163226 299512 163282 299568
rect 163410 299512 163466 299568
rect 56506 298016 56562 298072
rect 57886 298016 57942 298072
rect 59266 298016 59322 298072
rect 60646 298016 60702 298072
rect 62026 298016 62082 298072
rect 63406 298016 63462 298072
rect 64786 298016 64842 298072
rect 66166 298016 66222 298072
rect 67546 298016 67602 298072
rect 68742 298016 68798 298072
rect 70306 298016 70362 298072
rect 71686 298016 71742 298072
rect 73066 298016 73122 298072
rect 74446 298016 74502 298072
rect 75826 298016 75882 298072
rect 77022 298016 77078 298072
rect 78494 298016 78550 298072
rect 79966 298016 80022 298072
rect 80702 298016 80758 298072
rect 81254 298016 81310 298072
rect 82726 298016 82782 298072
rect 83370 298016 83426 298072
rect 84014 298016 84070 298072
rect 85486 298016 85542 298072
rect 86222 298016 86278 298072
rect 86774 298016 86830 298072
rect 88154 298016 88210 298072
rect 89626 298016 89682 298072
rect 91006 298016 91062 298072
rect 92386 298016 92442 298072
rect 93766 298016 93822 298072
rect 95146 298016 95202 298072
rect 96434 298016 96490 298072
rect 97906 298016 97962 298072
rect 99194 298016 99250 298072
rect 102046 298016 102102 298072
rect 106186 298016 106242 298072
rect 108486 298016 108542 298072
rect 111706 298016 111762 298072
rect 114466 298016 114522 298072
rect 115938 298016 115994 298072
rect 117410 298016 117466 298072
rect 121366 298016 121422 298072
rect 124126 298016 124182 298072
rect 125874 298016 125930 298072
rect 129646 298016 129702 298072
rect 133786 298016 133842 298072
rect 136086 298036 136142 298072
rect 136086 298016 136088 298036
rect 136088 298016 136140 298036
rect 136140 298016 136142 298036
rect 60554 297880 60610 297936
rect 66166 230016 66222 230072
rect 64786 229880 64842 229936
rect 68834 297900 68890 297936
rect 68834 297880 68836 297900
rect 68836 297880 68888 297900
rect 68888 297880 68890 297900
rect 68834 297744 68890 297800
rect 70306 239400 70362 239456
rect 74354 297880 74410 297936
rect 74354 230152 74410 230208
rect 77114 297880 77170 297936
rect 77206 297744 77262 297800
rect 78586 297880 78642 297936
rect 88246 297880 88302 297936
rect 90914 297880 90970 297936
rect 92294 297880 92350 297936
rect 93674 297880 93730 297936
rect 96526 297880 96582 297936
rect 99102 297880 99158 297936
rect 99286 297744 99342 297800
rect 104806 296792 104862 296848
rect 107658 223524 107660 223544
rect 107660 223524 107712 223544
rect 107712 223524 107714 223544
rect 107658 223488 107714 223524
rect 107658 217776 107714 217832
rect 107658 188808 107714 188864
rect 107658 186088 107714 186144
rect 107658 180648 107714 180704
rect 107658 177964 107660 177984
rect 107660 177964 107712 177984
rect 107712 177964 107714 177984
rect 107658 177928 107714 177964
rect 107658 172352 107714 172408
rect 107658 169668 107660 169688
rect 107660 169668 107712 169688
rect 107712 169668 107714 169688
rect 107658 169632 107714 169668
rect 108486 226208 108542 226264
rect 108578 215192 108634 215248
rect 108670 212472 108726 212528
rect 108762 206896 108818 206952
rect 108854 196832 108910 196888
rect 109406 209616 109462 209672
rect 139306 298016 139362 298072
rect 141054 298016 141110 298072
rect 146206 298016 146262 298072
rect 178682 379208 178738 379264
rect 178682 319368 178738 319424
rect 178958 317736 179014 317792
rect 178958 316376 179014 316432
rect 178590 314880 178646 314936
rect 178682 313656 178738 313712
rect 216678 336796 216734 336832
rect 216678 336776 216680 336796
rect 216680 336776 216732 336796
rect 216732 336776 216734 336796
rect 217322 335824 217378 335880
rect 216678 309848 216734 309904
rect 216770 308352 216826 308408
rect 217506 329840 217562 329896
rect 217966 333648 218022 333704
rect 217874 308352 217930 308408
rect 217874 307944 217930 308000
rect 251822 459856 251878 459912
rect 252098 461624 252154 461680
rect 376942 466792 376998 466848
rect 252466 466520 252522 466576
rect 376942 464208 376998 464264
rect 376942 461624 376998 461680
rect 376942 459040 376998 459096
rect 376942 456456 376998 456512
rect 376942 454008 376998 454064
rect 376850 451424 376906 451480
rect 376942 448840 376998 448896
rect 376942 446256 376998 446312
rect 376850 443672 376906 443728
rect 376942 441224 376998 441280
rect 248510 386280 248566 386336
rect 252558 386280 252614 386336
rect 255318 386280 255374 386336
rect 258262 386280 258318 386336
rect 260838 386280 260894 386336
rect 263598 386280 263654 386336
rect 264978 386280 265034 386336
rect 268106 386280 268162 386336
rect 270498 386280 270554 386336
rect 273258 386280 273314 386336
rect 249798 386008 249854 386064
rect 277950 386280 278006 386336
rect 280158 386280 280214 386336
rect 288438 386280 288494 386336
rect 285678 386144 285734 386200
rect 289818 386144 289874 386200
rect 295338 386280 295394 386336
rect 298098 385872 298154 385928
rect 304998 386280 305054 386336
rect 302238 385872 302294 385928
rect 310518 386280 310574 386336
rect 313278 386280 313334 386336
rect 317418 386280 317474 386336
rect 320178 386280 320234 386336
rect 322938 386280 322994 386336
rect 316038 386008 316094 386064
rect 338118 386280 338174 386336
rect 339498 386280 339554 386336
rect 276018 385056 276074 385112
rect 282918 385056 282974 385112
rect 292578 385056 292634 385112
rect 300858 385056 300914 385112
rect 307758 385056 307814 385112
rect 325882 385056 325938 385112
rect 350998 385056 351054 385112
rect 235998 298016 236054 298072
rect 238114 298016 238170 298072
rect 242806 298016 242862 298072
rect 247038 298016 247094 298072
rect 248418 298016 248474 298072
rect 249798 298016 249854 298072
rect 251086 298016 251142 298072
rect 251362 298016 251418 298072
rect 251546 298016 251602 298072
rect 252558 298016 252614 298072
rect 258170 298016 258226 298072
rect 259458 298016 259514 298072
rect 260194 298016 260250 298072
rect 261114 298016 261170 298072
rect 263690 298016 263746 298072
rect 265070 298016 265126 298072
rect 265346 298016 265402 298072
rect 266358 298016 266414 298072
rect 267830 298016 267886 298072
rect 269762 298016 269818 298072
rect 270498 298016 270554 298072
rect 271878 298016 271934 298072
rect 273258 298016 273314 298072
rect 274638 298016 274694 298072
rect 276018 298016 276074 298072
rect 276754 298016 276810 298072
rect 277490 298016 277546 298072
rect 278778 298016 278834 298072
rect 280158 298016 280214 298072
rect 282918 298016 282974 298072
rect 285954 298016 286010 298072
rect 287610 298016 287666 298072
rect 290002 298016 290058 298072
rect 292578 298016 292634 298072
rect 295338 298016 295394 298072
rect 298466 298016 298522 298072
rect 300858 298016 300914 298072
rect 302330 298016 302386 298072
rect 305090 298016 305146 298072
rect 308586 298016 308642 298072
rect 310978 298016 311034 298072
rect 313278 298016 313334 298072
rect 315762 298016 315818 298072
rect 317418 298016 317474 298072
rect 320914 298016 320970 298072
rect 322938 298016 322994 298072
rect 325698 298016 325754 298072
rect 343178 298036 343234 298072
rect 343178 298016 343180 298036
rect 343180 298016 343232 298036
rect 343232 298016 343234 298036
rect 237286 297880 237342 297936
rect 240046 296792 240102 296848
rect 248326 297880 248382 297936
rect 256606 296928 256662 296984
rect 255318 296792 255374 296848
rect 256698 296792 256754 296848
rect 258078 296792 258134 296848
rect 258354 297744 258410 297800
rect 258354 295976 258410 296032
rect 259366 229472 259422 229528
rect 110326 228928 110382 228984
rect 109590 220428 109646 220484
rect 109498 204856 109554 204912
rect 109314 202272 109370 202328
rect 109222 199552 109278 199608
rect 109130 194112 109186 194168
rect 260930 296792 260986 296848
rect 263598 297880 263654 297936
rect 262218 296792 262274 296848
rect 259918 227976 259974 228032
rect 259826 226208 259882 226264
rect 259734 209072 259790 209128
rect 259642 205536 259698 205592
rect 259550 202680 259606 202736
rect 259458 191528 259514 191584
rect 109038 191392 109094 191448
rect 108946 183368 109002 183424
rect 108394 175208 108450 175264
rect 108210 166912 108266 166968
rect 107658 164056 107714 164112
rect 260286 198804 260342 198860
rect 260194 192548 260250 192604
rect 260102 187652 260158 187708
rect 260010 172352 260066 172408
rect 261206 212200 261262 212256
rect 262218 189932 262220 189952
rect 262220 189932 262272 189952
rect 262272 189932 262274 189952
rect 262218 189896 262274 189932
rect 262678 220224 262734 220280
rect 262954 223080 263010 223136
rect 262862 221720 262918 221776
rect 262678 215192 262734 215248
rect 262586 206896 262642 206952
rect 262494 201048 262550 201104
rect 262402 195880 262458 195936
rect 262310 182008 262366 182064
rect 261114 180240 261170 180296
rect 261022 178744 261078 178800
rect 260930 173848 260986 173904
rect 260838 169224 260894 169280
rect 259918 165280 259974 165336
rect 259826 162696 259882 162752
rect 107658 161372 107660 161392
rect 107660 161372 107712 161392
rect 107712 161372 107714 161392
rect 107658 161336 107714 161372
rect 263506 224576 263562 224632
rect 263506 217948 263508 217968
rect 263508 217948 263560 217968
rect 263560 217948 263562 217968
rect 263506 217912 263562 217948
rect 263506 216416 263562 216472
rect 263506 213560 263562 213616
rect 263506 210568 263562 210624
rect 263506 203904 263562 203960
rect 263046 161064 263102 161120
rect 216770 160384 216826 160440
rect 218886 160384 218942 160440
rect 215850 158480 215906 158536
rect 220726 158344 220782 158400
rect 223670 158208 223726 158264
rect 222290 158072 222346 158128
rect 228914 158072 228970 158128
rect 258170 158208 258226 158264
rect 251914 157936 251970 157992
rect 266450 297880 266506 297936
rect 268014 297880 268070 297936
rect 270590 297880 270646 297936
rect 273350 297880 273406 297936
rect 273442 297744 273498 297800
rect 276662 296928 276718 296984
rect 343362 298052 343364 298072
rect 343364 298052 343416 298072
rect 343416 298052 343418 298072
rect 343362 298016 343418 298052
rect 256698 119448 256754 119504
rect 342258 119448 342314 119504
rect 256698 118652 256754 118688
rect 256698 118632 256700 118652
rect 256700 118632 256752 118652
rect 256752 118632 256754 118652
rect 342258 118632 342314 118688
rect 256790 117816 256846 117872
rect 342350 117816 342406 117872
rect 256698 117000 256754 117056
rect 342258 117000 342314 117056
rect 256790 116184 256846 116240
rect 342350 116184 342406 116240
rect 256698 115368 256754 115424
rect 342258 115368 342314 115424
rect 256790 114552 256846 114608
rect 342350 114552 342406 114608
rect 256698 113736 256754 113792
rect 342258 113736 342314 113792
rect 256698 113076 256754 113112
rect 342258 113092 342260 113112
rect 342260 113092 342312 113112
rect 342312 113092 342314 113112
rect 256698 113056 256700 113076
rect 256700 113056 256752 113076
rect 256752 113056 256754 113076
rect 342258 113056 342314 113092
rect 256790 112240 256846 112296
rect 342350 112240 342406 112296
rect 256698 111424 256754 111480
rect 342258 111424 342314 111480
rect 256790 110608 256846 110664
rect 342350 110608 342406 110664
rect 256698 109792 256754 109848
rect 342258 109792 342314 109848
rect 256698 108976 256754 109032
rect 342258 108996 342314 109032
rect 342258 108976 342260 108996
rect 342260 108976 342312 108996
rect 342312 108976 342314 108996
rect 256790 108160 256846 108216
rect 342350 108160 342406 108216
rect 256698 107344 256754 107400
rect 342258 107344 342314 107400
rect 256790 106664 256846 106720
rect 342350 106664 342406 106720
rect 256698 105848 256754 105904
rect 342258 105848 342314 105904
rect 256790 105032 256846 105088
rect 342350 105032 342406 105088
rect 256698 104216 256754 104272
rect 342258 104216 342314 104272
rect 256698 103420 256754 103456
rect 342258 103436 342260 103456
rect 342260 103436 342312 103456
rect 342312 103436 342314 103456
rect 256698 103400 256700 103420
rect 256700 103400 256752 103420
rect 256752 103400 256754 103420
rect 342258 103400 342314 103436
rect 256790 102584 256846 102640
rect 342350 102584 342406 102640
rect 256698 101768 256754 101824
rect 342258 101768 342314 101824
rect 256790 100952 256846 101008
rect 342350 100952 342406 101008
rect 256698 100272 256754 100328
rect 342258 100272 342314 100328
rect 256790 99456 256846 99512
rect 342350 99456 342406 99512
rect 256698 98640 256754 98696
rect 342258 98640 342314 98696
rect 256698 97860 256700 97880
rect 256700 97860 256752 97880
rect 256752 97860 256754 97880
rect 256698 97824 256754 97860
rect 342258 97824 342314 97880
rect 256790 97008 256846 97064
rect 342350 97008 342406 97064
rect 256698 96192 256754 96248
rect 342258 96192 342314 96248
rect 256790 95376 256846 95432
rect 342350 95376 342406 95432
rect 256698 94560 256754 94616
rect 342258 94560 342314 94616
rect 256698 93764 256754 93800
rect 342258 93780 342260 93800
rect 342260 93780 342312 93800
rect 342312 93780 342314 93800
rect 256698 93744 256700 93764
rect 256700 93744 256752 93764
rect 256752 93744 256754 93764
rect 342258 93744 342314 93780
rect 256790 93064 256846 93120
rect 342350 93064 342406 93120
rect 256698 92248 256754 92304
rect 342258 92248 342314 92304
rect 256790 91432 256846 91488
rect 342350 91432 342406 91488
rect 256698 90616 256754 90672
rect 342258 90616 342314 90672
rect 256790 89800 256846 89856
rect 342350 89800 342406 89856
rect 256698 88984 256754 89040
rect 342258 88984 342314 89040
rect 256698 88204 256700 88224
rect 256700 88204 256752 88224
rect 256752 88204 256754 88224
rect 256698 88168 256754 88204
rect 342258 88168 342314 88224
rect 256790 87352 256846 87408
rect 342350 87352 342406 87408
rect 256698 86672 256754 86728
rect 342258 86672 342314 86728
rect 256790 85856 256846 85912
rect 342350 85856 342406 85912
rect 256698 85040 256754 85096
rect 342258 85040 342314 85096
rect 256790 84224 256846 84280
rect 342350 84224 342406 84280
rect 256698 83408 256754 83464
rect 342258 83408 342314 83464
rect 256698 82592 256754 82648
rect 342258 82592 342314 82648
rect 256790 81776 256846 81832
rect 342350 81776 342406 81832
rect 256698 80960 256754 81016
rect 342258 80960 342314 81016
rect 256790 80280 256846 80336
rect 342350 80280 342406 80336
rect 256698 79464 256754 79520
rect 342258 79464 342314 79520
rect 256790 78648 256846 78704
rect 342350 78648 342406 78704
rect 256698 77832 256754 77888
rect 342258 77832 342314 77888
rect 256698 77016 256754 77072
rect 342258 77016 342314 77072
rect 256790 76200 256846 76256
rect 342350 76200 342406 76256
rect 256698 75384 256754 75440
rect 342258 75384 342314 75440
rect 256790 74568 256846 74624
rect 342350 74568 342406 74624
rect 256698 73752 256754 73808
rect 342258 73752 342314 73808
rect 256698 73092 256754 73128
rect 342258 73108 342260 73128
rect 342260 73108 342312 73128
rect 342312 73108 342314 73128
rect 256698 73072 256700 73092
rect 256700 73072 256752 73092
rect 256752 73072 256754 73092
rect 342258 73072 342314 73108
rect 256790 72256 256846 72312
rect 342350 72256 342406 72312
rect 256698 71440 256754 71496
rect 342258 71440 342314 71496
rect 256790 70624 256846 70680
rect 342350 70624 342406 70680
rect 256698 69808 256754 69864
rect 342258 69808 342314 69864
rect 256790 68992 256846 69048
rect 342350 68992 342406 69048
rect 256698 68176 256754 68232
rect 342258 68176 342314 68232
rect 256698 67360 256754 67416
rect 342258 67360 342314 67416
rect 256790 66680 256846 66736
rect 342350 66680 342406 66736
rect 256698 65864 256754 65920
rect 342258 65864 342314 65920
rect 256790 65048 256846 65104
rect 342350 65048 342406 65104
rect 256698 64232 256754 64288
rect 342258 64232 342314 64288
rect 256698 63436 256754 63472
rect 342258 63452 342260 63472
rect 342260 63452 342312 63472
rect 342312 63452 342314 63472
rect 256698 63416 256700 63436
rect 256700 63416 256752 63436
rect 256752 63416 256754 63436
rect 342258 63416 342314 63452
rect 256790 62600 256846 62656
rect 342350 62600 342406 62656
rect 256698 61784 256754 61840
rect 342258 61784 342314 61840
rect 256790 60968 256846 61024
rect 342350 60968 342406 61024
rect 256698 60288 256754 60344
rect 342258 60288 342314 60344
rect 256790 59472 256846 59528
rect 342350 59472 342406 59528
rect 256698 58656 256754 58712
rect 342258 58656 342314 58712
rect 256698 57860 256754 57896
rect 342258 57876 342260 57896
rect 342260 57876 342312 57896
rect 342312 57876 342314 57896
rect 256698 57840 256700 57860
rect 256700 57840 256752 57860
rect 256752 57840 256754 57860
rect 342258 57840 342314 57876
rect 256790 57024 256846 57080
rect 342350 57024 342406 57080
rect 256698 56208 256754 56264
rect 342258 56208 342314 56264
rect 256790 55392 256846 55448
rect 342350 55392 342406 55448
rect 256698 54576 256754 54632
rect 342258 54576 342314 54632
rect 256698 53760 256754 53816
rect 342258 53780 342314 53816
rect 342258 53760 342260 53780
rect 342260 53760 342312 53780
rect 342312 53760 342314 53780
rect 256790 53080 256846 53136
rect 342350 53080 342406 53136
rect 256698 52300 256700 52320
rect 256700 52300 256752 52320
rect 256752 52300 256754 52320
rect 256698 52264 256754 52300
rect 342258 52264 342314 52320
rect 256790 51448 256846 51504
rect 342350 51448 342406 51504
rect 256698 50632 256754 50688
rect 342258 50632 342314 50688
rect 256790 49816 256846 49872
rect 342350 49816 342406 49872
rect 256698 49000 256754 49056
rect 342258 49000 342314 49056
rect 256698 48204 256754 48240
rect 342258 48220 342260 48240
rect 342260 48220 342312 48240
rect 342312 48220 342314 48240
rect 256698 48184 256700 48204
rect 256700 48184 256752 48204
rect 256752 48184 256754 48204
rect 342258 48184 342314 48220
rect 256790 47368 256846 47424
rect 342350 47368 342406 47424
rect 256698 46688 256754 46744
rect 359278 379344 359334 379400
rect 359186 319912 359242 319968
rect 359094 318280 359150 318336
rect 359002 316920 359058 316976
rect 358910 315424 358966 315480
rect 358818 314200 358874 314256
rect 342258 46688 342314 46744
rect 256790 45872 256846 45928
rect 342350 45872 342406 45928
rect 256698 45056 256754 45112
rect 342258 45056 342314 45112
rect 256790 44240 256846 44296
rect 342350 44240 342406 44296
rect 256698 43424 256754 43480
rect 342258 43424 342314 43480
rect 256698 42644 256700 42664
rect 256700 42644 256752 42664
rect 256752 42644 256754 42664
rect 256698 42608 256754 42644
rect 342258 42608 342314 42664
rect 256790 41792 256846 41848
rect 342350 41792 342406 41848
rect 256698 40976 256754 41032
rect 579894 537784 579950 537840
rect 580170 524456 580226 524512
rect 580262 484608 580318 484664
rect 580170 471416 580226 471472
rect 579802 431568 579858 431624
rect 580170 418240 580226 418296
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 342258 40976 342314 41032
rect 256790 40296 256846 40352
rect 342350 40296 342406 40352
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 579852 480 580092
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect 376937 548722 377003 548725
rect 376937 548720 380052 548722
rect 376937 548664 376942 548720
rect 376998 548664 380052 548720
rect 376937 548662 380052 548664
rect 376937 548659 377003 548662
rect 376937 546138 377003 546141
rect 376937 546136 380052 546138
rect 376937 546080 376942 546136
rect 376998 546080 380052 546136
rect 376937 546078 380052 546080
rect 376937 546075 377003 546078
rect 376845 543554 376911 543557
rect 376845 543552 380052 543554
rect 376845 543496 376850 543552
rect 376906 543496 380052 543552
rect 376845 543494 380052 543496
rect 376845 543491 376911 543494
rect 377397 540970 377463 540973
rect 377397 540968 380052 540970
rect -960 540684 480 540924
rect 377397 540912 377402 540968
rect 377458 540912 380052 540968
rect 377397 540910 380052 540912
rect 377397 540907 377463 540910
rect 376937 538386 377003 538389
rect 376937 538384 380052 538386
rect 376937 538328 376942 538384
rect 376998 538328 380052 538384
rect 376937 538326 380052 538328
rect 376937 538323 377003 538326
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 376937 535938 377003 535941
rect 376937 535936 380052 535938
rect 376937 535880 376942 535936
rect 376998 535880 380052 535936
rect 376937 535878 380052 535880
rect 376937 535875 377003 535878
rect 376937 533354 377003 533357
rect 376937 533352 380052 533354
rect 376937 533296 376942 533352
rect 376998 533296 380052 533352
rect 376937 533294 380052 533296
rect 376937 533291 377003 533294
rect 377489 530770 377555 530773
rect 377489 530768 380052 530770
rect 377489 530712 377494 530768
rect 377550 530712 380052 530768
rect 377489 530710 380052 530712
rect 377489 530707 377555 530710
rect 376937 528186 377003 528189
rect 376937 528184 380052 528186
rect 376937 528128 376942 528184
rect 376998 528128 380052 528184
rect 376937 528126 380052 528128
rect 376937 528123 377003 528126
rect -960 527764 480 528004
rect 376937 525602 377003 525605
rect 376937 525600 380052 525602
rect 376937 525544 376942 525600
rect 376998 525544 380052 525600
rect 376937 525542 380052 525544
rect 376937 525539 377003 525542
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 376937 523154 377003 523157
rect 376937 523152 380052 523154
rect 376937 523096 376942 523152
rect 376998 523096 380052 523152
rect 376937 523094 380052 523096
rect 376937 523091 377003 523094
rect 377581 520570 377647 520573
rect 377581 520568 380052 520570
rect 377581 520512 377586 520568
rect 377642 520512 380052 520568
rect 377581 520510 380052 520512
rect 377581 520507 377647 520510
rect 376937 517986 377003 517989
rect 376937 517984 380052 517986
rect 376937 517928 376942 517984
rect 376998 517928 380052 517984
rect 376937 517926 380052 517928
rect 376937 517923 377003 517926
rect 376937 515402 377003 515405
rect 376937 515400 380052 515402
rect 376937 515344 376942 515400
rect 376998 515344 380052 515400
rect 376937 515342 380052 515344
rect 376937 515339 377003 515342
rect -960 514708 480 514948
rect 376937 512818 377003 512821
rect 376937 512816 380052 512818
rect 376937 512760 376942 512816
rect 376998 512760 380052 512816
rect 376937 512758 380052 512760
rect 376937 512755 377003 512758
rect 583520 511172 584960 511412
rect 376937 510234 377003 510237
rect 376937 510232 380052 510234
rect 376937 510176 376942 510232
rect 376998 510176 380052 510232
rect 376937 510174 380052 510176
rect 376937 510171 377003 510174
rect 377673 507786 377739 507789
rect 377673 507784 380052 507786
rect 377673 507728 377678 507784
rect 377734 507728 380052 507784
rect 377673 507726 380052 507728
rect 377673 507723 377739 507726
rect 377765 505202 377831 505205
rect 377765 505200 380052 505202
rect 377765 505144 377770 505200
rect 377826 505144 380052 505200
rect 377765 505142 380052 505144
rect 377765 505139 377831 505142
rect 377857 502618 377923 502621
rect 377857 502616 380052 502618
rect 377857 502560 377862 502616
rect 377918 502560 380052 502616
rect 377857 502558 380052 502560
rect 377857 502555 377923 502558
rect -960 501652 480 501892
rect 377949 500034 378015 500037
rect 377949 500032 380052 500034
rect 377949 499976 377954 500032
rect 378010 499976 380052 500032
rect 377949 499974 380052 499976
rect 377949 499971 378015 499974
rect 249934 499354 249994 499460
rect 252461 499354 252527 499357
rect 249934 499352 252527 499354
rect 249934 499296 252466 499352
rect 252522 499296 252527 499352
rect 249934 499294 252527 499296
rect 252461 499291 252527 499294
rect 251817 499082 251883 499085
rect 249934 499080 251883 499082
rect 249934 499024 251822 499080
rect 251878 499024 251883 499080
rect 249934 499022 251883 499024
rect 249934 498508 249994 499022
rect 251817 499019 251883 499022
rect 252461 497858 252527 497861
rect 249934 497856 252527 497858
rect 249934 497800 252466 497856
rect 252522 497800 252527 497856
rect 583520 497844 584960 498084
rect 249934 497798 252527 497800
rect 249934 497556 249994 497798
rect 252461 497795 252527 497798
rect 378041 497450 378107 497453
rect 378041 497448 380052 497450
rect 378041 497392 378046 497448
rect 378102 497392 380052 497448
rect 378041 497390 380052 497392
rect 378041 497387 378107 497390
rect 252461 496770 252527 496773
rect 249934 496768 252527 496770
rect 249934 496712 252466 496768
rect 252522 496712 252527 496768
rect 249934 496710 252527 496712
rect 249934 496604 249994 496710
rect 252461 496707 252527 496710
rect 252369 496226 252435 496229
rect 249934 496224 252435 496226
rect 249934 496168 252374 496224
rect 252430 496168 252435 496224
rect 249934 496166 252435 496168
rect 249934 495652 249994 496166
rect 252369 496163 252435 496166
rect 251909 495274 251975 495277
rect 249934 495272 251975 495274
rect 249934 495216 251914 495272
rect 251970 495216 251975 495272
rect 249934 495214 251975 495216
rect 249934 494700 249994 495214
rect 251909 495211 251975 495214
rect 377397 495002 377463 495005
rect 377397 495000 380052 495002
rect 377397 494944 377402 495000
rect 377458 494944 380052 495000
rect 377397 494942 380052 494944
rect 377397 494939 377463 494942
rect 252461 494050 252527 494053
rect 249934 494048 252527 494050
rect 249934 493992 252466 494048
rect 252522 493992 252527 494048
rect 249934 493990 252527 493992
rect 249934 493884 249994 493990
rect 252461 493987 252527 493990
rect 252369 493506 252435 493509
rect 249934 493504 252435 493506
rect 249934 493448 252374 493504
rect 252430 493448 252435 493504
rect 249934 493446 252435 493448
rect 249934 492932 249994 493446
rect 252369 493443 252435 493446
rect 376937 492418 377003 492421
rect 376937 492416 380052 492418
rect 376937 492360 376942 492416
rect 376998 492360 380052 492416
rect 376937 492358 380052 492360
rect 376937 492355 377003 492358
rect 252461 492146 252527 492149
rect 249934 492144 252527 492146
rect 249934 492088 252466 492144
rect 252522 492088 252527 492144
rect 249934 492086 252527 492088
rect 249934 491980 249994 492086
rect 252461 492083 252527 492086
rect 252001 491194 252067 491197
rect 249934 491192 252067 491194
rect 249934 491136 252006 491192
rect 252062 491136 252067 491192
rect 249934 491134 252067 491136
rect 249934 491028 249994 491134
rect 252001 491131 252067 491134
rect 251909 490650 251975 490653
rect 249934 490648 251975 490650
rect 249934 490592 251914 490648
rect 251970 490592 251975 490648
rect 249934 490590 251975 490592
rect 249934 490076 249994 490590
rect 251909 490587 251975 490590
rect 376937 489834 377003 489837
rect 376937 489832 380052 489834
rect 376937 489776 376942 489832
rect 376998 489776 380052 489832
rect 376937 489774 380052 489776
rect 376937 489771 377003 489774
rect 252461 489562 252527 489565
rect 249934 489560 252527 489562
rect 249934 489504 252466 489560
rect 252522 489504 252527 489560
rect 249934 489502 252527 489504
rect 249934 489124 249994 489502
rect 252461 489499 252527 489502
rect -960 488596 480 488836
rect 252461 488474 252527 488477
rect 249934 488472 252527 488474
rect 249934 488416 252466 488472
rect 252522 488416 252527 488472
rect 249934 488414 252527 488416
rect 249934 488308 249994 488414
rect 252461 488411 252527 488414
rect 252093 487930 252159 487933
rect 249934 487928 252159 487930
rect 249934 487872 252098 487928
rect 252154 487872 252159 487928
rect 249934 487870 252159 487872
rect 249934 487356 249994 487870
rect 252093 487867 252159 487870
rect 376937 487250 377003 487253
rect 376937 487248 380052 487250
rect 376937 487192 376942 487248
rect 376998 487192 380052 487248
rect 376937 487190 380052 487192
rect 376937 487187 377003 487190
rect 251265 486978 251331 486981
rect 249934 486976 251331 486978
rect 249934 486920 251270 486976
rect 251326 486920 251331 486976
rect 249934 486918 251331 486920
rect 249934 486404 249994 486918
rect 251265 486915 251331 486918
rect 251357 485618 251423 485621
rect 249934 485616 251423 485618
rect 249934 485560 251362 485616
rect 251418 485560 251423 485616
rect 249934 485558 251423 485560
rect 249934 485452 249994 485558
rect 251357 485555 251423 485558
rect 251725 485074 251791 485077
rect 249934 485072 251791 485074
rect 249934 485016 251730 485072
rect 251786 485016 251791 485072
rect 249934 485014 251791 485016
rect 249934 484500 249994 485014
rect 251725 485011 251791 485014
rect 377489 484666 377555 484669
rect 580257 484666 580323 484669
rect 583520 484666 584960 484756
rect 377489 484664 380052 484666
rect 377489 484608 377494 484664
rect 377550 484608 380052 484664
rect 377489 484606 380052 484608
rect 580257 484664 584960 484666
rect 580257 484608 580262 484664
rect 580318 484608 584960 484664
rect 580257 484606 584960 484608
rect 377489 484603 377555 484606
rect 580257 484603 580323 484606
rect 583520 484516 584960 484606
rect 251725 483986 251791 483989
rect 249934 483984 251791 483986
rect 249934 483928 251730 483984
rect 251786 483928 251791 483984
rect 249934 483926 251791 483928
rect 249934 483548 249994 483926
rect 251725 483923 251791 483926
rect 252461 482898 252527 482901
rect 249934 482896 252527 482898
rect 249934 482840 252466 482896
rect 252522 482840 252527 482896
rect 249934 482838 252527 482840
rect 249934 482732 249994 482838
rect 252461 482835 252527 482838
rect 252369 482354 252435 482357
rect 249934 482352 252435 482354
rect 249934 482296 252374 482352
rect 252430 482296 252435 482352
rect 249934 482294 252435 482296
rect 249934 481780 249994 482294
rect 252369 482291 252435 482294
rect 377213 482218 377279 482221
rect 377213 482216 380052 482218
rect 377213 482160 377218 482216
rect 377274 482160 380052 482216
rect 377213 482158 380052 482160
rect 377213 482155 377279 482158
rect 251725 481266 251791 481269
rect 249934 481264 251791 481266
rect 249934 481208 251730 481264
rect 251786 481208 251791 481264
rect 249934 481206 251791 481208
rect 249934 480828 249994 481206
rect 251725 481203 251791 481206
rect 252461 480042 252527 480045
rect 249934 480040 252527 480042
rect 249934 479984 252466 480040
rect 252522 479984 252527 480040
rect 249934 479982 252527 479984
rect 249934 479876 249994 479982
rect 252461 479979 252527 479982
rect 377029 479634 377095 479637
rect 377029 479632 380052 479634
rect 377029 479576 377034 479632
rect 377090 479576 380052 479632
rect 377029 479574 380052 479576
rect 377029 479571 377095 479574
rect 251817 479498 251883 479501
rect 249934 479496 251883 479498
rect 249934 479440 251822 479496
rect 251878 479440 251883 479496
rect 249934 479438 251883 479440
rect 249934 478924 249994 479438
rect 251817 479435 251883 479438
rect 252001 478546 252067 478549
rect 249934 478544 252067 478546
rect 249934 478488 252006 478544
rect 252062 478488 252067 478544
rect 249934 478486 252067 478488
rect 249934 477972 249994 478486
rect 252001 478483 252067 478486
rect 251909 477458 251975 477461
rect 249934 477456 251975 477458
rect 249934 477400 251914 477456
rect 251970 477400 251975 477456
rect 249934 477398 251975 477400
rect 249934 477156 249994 477398
rect 251909 477395 251975 477398
rect 376937 477050 377003 477053
rect 376937 477048 380052 477050
rect 376937 476992 376942 477048
rect 376998 476992 380052 477048
rect 376937 476990 380052 476992
rect 376937 476987 377003 476990
rect 251725 476778 251791 476781
rect 249934 476776 251791 476778
rect 249934 476720 251730 476776
rect 251786 476720 251791 476776
rect 249934 476718 251791 476720
rect 249934 476204 249994 476718
rect 251725 476715 251791 476718
rect -960 475540 480 475780
rect 252461 475690 252527 475693
rect 249934 475688 252527 475690
rect 249934 475632 252466 475688
rect 252522 475632 252527 475688
rect 249934 475630 252527 475632
rect 249934 475252 249994 475630
rect 252461 475627 252527 475630
rect 252461 474466 252527 474469
rect 249934 474464 252527 474466
rect 249934 474408 252466 474464
rect 252522 474408 252527 474464
rect 249934 474406 252527 474408
rect 249934 474300 249994 474406
rect 252461 474403 252527 474406
rect 376937 474466 377003 474469
rect 376937 474464 380052 474466
rect 376937 474408 376942 474464
rect 376998 474408 380052 474464
rect 376937 474406 380052 474408
rect 376937 474403 377003 474406
rect 251909 473922 251975 473925
rect 249934 473920 251975 473922
rect 249934 473864 251914 473920
rect 251970 473864 251975 473920
rect 249934 473862 251975 473864
rect 249934 473348 249994 473862
rect 251909 473859 251975 473862
rect 251541 472970 251607 472973
rect 249934 472968 251607 472970
rect 249934 472912 251546 472968
rect 251602 472912 251607 472968
rect 249934 472910 251607 472912
rect 249934 472396 249994 472910
rect 251541 472907 251607 472910
rect 376937 471882 377003 471885
rect 376937 471880 380052 471882
rect 376937 471824 376942 471880
rect 376998 471824 380052 471880
rect 376937 471822 380052 471824
rect 376937 471819 377003 471822
rect 249934 471474 249994 471580
rect 252461 471474 252527 471477
rect 249934 471472 252527 471474
rect 249934 471416 252466 471472
rect 252522 471416 252527 471472
rect 249934 471414 252527 471416
rect 252461 471411 252527 471414
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 252461 470794 252527 470797
rect 249934 470792 252527 470794
rect 249934 470736 252466 470792
rect 252522 470736 252527 470792
rect 249934 470734 252527 470736
rect 249934 470628 249994 470734
rect 252461 470731 252527 470734
rect 249934 469298 249994 469676
rect 252461 469298 252527 469301
rect 249934 469296 252527 469298
rect 249934 469240 252466 469296
rect 252522 469240 252527 469296
rect 249934 469238 252527 469240
rect 252461 469235 252527 469238
rect 376937 469298 377003 469301
rect 376937 469296 380052 469298
rect 376937 469240 376942 469296
rect 376998 469240 380052 469296
rect 376937 469238 380052 469240
rect 376937 469235 377003 469238
rect 249934 468210 249994 468724
rect 252369 468210 252435 468213
rect 249934 468208 252435 468210
rect 249934 468152 252374 468208
rect 252430 468152 252435 468208
rect 249934 468150 252435 468152
rect 252369 468147 252435 468150
rect 249934 467258 249994 467772
rect 251541 467258 251607 467261
rect 249934 467256 251607 467258
rect 249934 467200 251546 467256
rect 251602 467200 251607 467256
rect 249934 467198 251607 467200
rect 251541 467195 251607 467198
rect 376937 466850 377003 466853
rect 376937 466848 380052 466850
rect 249934 466578 249994 466820
rect 376937 466792 376942 466848
rect 376998 466792 380052 466848
rect 376937 466790 380052 466792
rect 376937 466787 377003 466790
rect 252461 466578 252527 466581
rect 249934 466576 252527 466578
rect 249934 466520 252466 466576
rect 252522 466520 252527 466576
rect 249934 466518 252527 466520
rect 252461 466515 252527 466518
rect 249934 465490 249994 466004
rect 252277 465490 252343 465493
rect 249934 465488 252343 465490
rect 249934 465432 252282 465488
rect 252338 465432 252343 465488
rect 249934 465430 252343 465432
rect 252277 465427 252343 465430
rect 249934 464538 249994 465052
rect 251265 464538 251331 464541
rect 249934 464536 251331 464538
rect 249934 464480 251270 464536
rect 251326 464480 251331 464536
rect 249934 464478 251331 464480
rect 251265 464475 251331 464478
rect 376937 464266 377003 464269
rect 376937 464264 380052 464266
rect 376937 464208 376942 464264
rect 376998 464208 380052 464264
rect 376937 464206 380052 464208
rect 376937 464203 377003 464206
rect 249934 463722 249994 464100
rect 252185 463722 252251 463725
rect 249934 463720 252251 463722
rect 249934 463664 252190 463720
rect 252246 463664 252251 463720
rect 249934 463662 252251 463664
rect 252185 463659 252251 463662
rect -960 462484 480 462724
rect 249934 462634 249994 463148
rect 252001 462634 252067 462637
rect 249934 462632 252067 462634
rect 249934 462576 252006 462632
rect 252062 462576 252067 462632
rect 249934 462574 252067 462576
rect 252001 462571 252067 462574
rect 249934 461682 249994 462196
rect 252093 461682 252159 461685
rect 249934 461680 252159 461682
rect 249934 461624 252098 461680
rect 252154 461624 252159 461680
rect 249934 461622 252159 461624
rect 252093 461619 252159 461622
rect 376937 461682 377003 461685
rect 376937 461680 380052 461682
rect 376937 461624 376942 461680
rect 376998 461624 380052 461680
rect 376937 461622 380052 461624
rect 376937 461619 377003 461622
rect 249934 461138 249994 461244
rect 251909 461138 251975 461141
rect 249934 461136 251975 461138
rect 249934 461080 251914 461136
rect 251970 461080 251975 461136
rect 249934 461078 251975 461080
rect 251909 461075 251975 461078
rect 249934 459914 249994 460428
rect 251817 459914 251883 459917
rect 249934 459912 251883 459914
rect 249934 459856 251822 459912
rect 251878 459856 251883 459912
rect 249934 459854 251883 459856
rect 251817 459851 251883 459854
rect 376937 459098 377003 459101
rect 376937 459096 380052 459098
rect 376937 459040 376942 459096
rect 376998 459040 380052 459096
rect 376937 459038 380052 459040
rect 376937 459035 377003 459038
rect 583520 457996 584960 458236
rect 376937 456514 377003 456517
rect 376937 456512 380052 456514
rect 376937 456456 376942 456512
rect 376998 456456 380052 456512
rect 376937 456454 380052 456456
rect 376937 456451 377003 456454
rect 376937 454066 377003 454069
rect 376937 454064 380052 454066
rect 376937 454008 376942 454064
rect 376998 454008 380052 454064
rect 376937 454006 380052 454008
rect 376937 454003 377003 454006
rect 376845 451482 376911 451485
rect 376845 451480 380052 451482
rect 376845 451424 376850 451480
rect 376906 451424 380052 451480
rect 376845 451422 380052 451424
rect 376845 451419 376911 451422
rect -960 449428 480 449668
rect 376937 448898 377003 448901
rect 376937 448896 380052 448898
rect 376937 448840 376942 448896
rect 376998 448840 380052 448896
rect 376937 448838 380052 448840
rect 376937 448835 377003 448838
rect 376937 446314 377003 446317
rect 376937 446312 380052 446314
rect 376937 446256 376942 446312
rect 376998 446256 380052 446312
rect 376937 446254 380052 446256
rect 376937 446251 377003 446254
rect 583520 444668 584960 444908
rect 376845 443730 376911 443733
rect 376845 443728 380052 443730
rect 376845 443672 376850 443728
rect 376906 443672 380052 443728
rect 376845 443670 380052 443672
rect 376845 443667 376911 443670
rect 376937 441282 377003 441285
rect 376937 441280 380052 441282
rect 376937 441224 376942 441280
rect 376998 441224 380052 441280
rect 376937 441222 380052 441224
rect 376937 441219 377003 441222
rect -960 436508 480 436748
rect 579797 431626 579863 431629
rect 583520 431626 584960 431716
rect 579797 431624 584960 431626
rect 579797 431568 579802 431624
rect 579858 431568 584960 431624
rect 579797 431566 584960 431568
rect 579797 431563 579863 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect 68737 386340 68803 386341
rect 68686 386338 68692 386340
rect 68646 386278 68692 386338
rect 68756 386336 68803 386340
rect 68798 386280 68803 386336
rect 68686 386276 68692 386278
rect 68756 386276 68803 386280
rect 71078 386276 71084 386340
rect 71148 386338 71154 386340
rect 71313 386338 71379 386341
rect 78489 386340 78555 386341
rect 78438 386338 78444 386340
rect 71148 386336 71379 386338
rect 71148 386280 71318 386336
rect 71374 386280 71379 386336
rect 71148 386278 71379 386280
rect 78398 386278 78444 386338
rect 78508 386336 78555 386340
rect 78550 386280 78555 386336
rect 71148 386276 71154 386278
rect 68737 386275 68803 386276
rect 71313 386275 71379 386278
rect 78438 386276 78444 386278
rect 78508 386276 78555 386280
rect 88558 386276 88564 386340
rect 88628 386338 88634 386340
rect 89161 386338 89227 386341
rect 88628 386336 89227 386338
rect 88628 386280 89166 386336
rect 89222 386280 89227 386336
rect 88628 386278 89227 386280
rect 88628 386276 88634 386278
rect 78489 386275 78555 386276
rect 89161 386275 89227 386278
rect 93526 386276 93532 386340
rect 93596 386338 93602 386340
rect 93761 386338 93827 386341
rect 93596 386336 93827 386338
rect 93596 386280 93766 386336
rect 93822 386280 93827 386336
rect 93596 386278 93827 386280
rect 93596 386276 93602 386278
rect 93761 386275 93827 386278
rect 96286 386276 96292 386340
rect 96356 386338 96362 386340
rect 96521 386338 96587 386341
rect 96356 386336 96587 386338
rect 96356 386280 96526 386336
rect 96582 386280 96587 386336
rect 96356 386278 96587 386280
rect 96356 386276 96362 386278
rect 96521 386275 96587 386278
rect 98494 386276 98500 386340
rect 98564 386338 98570 386340
rect 99281 386338 99347 386341
rect 98564 386336 99347 386338
rect 98564 386280 99286 386336
rect 99342 386280 99347 386336
rect 98564 386278 99347 386280
rect 98564 386276 98570 386278
rect 99281 386275 99347 386278
rect 100886 386276 100892 386340
rect 100956 386338 100962 386340
rect 102041 386338 102107 386341
rect 100956 386336 102107 386338
rect 100956 386280 102046 386336
rect 102102 386280 102107 386336
rect 100956 386278 102107 386280
rect 100956 386276 100962 386278
rect 102041 386275 102107 386278
rect 106038 386276 106044 386340
rect 106108 386338 106114 386340
rect 106181 386338 106247 386341
rect 106108 386336 106247 386338
rect 106108 386280 106186 386336
rect 106242 386280 106247 386336
rect 106108 386278 106247 386280
rect 106108 386276 106114 386278
rect 106181 386275 106247 386278
rect 108614 386276 108620 386340
rect 108684 386338 108690 386340
rect 108941 386338 109007 386341
rect 108684 386336 109007 386338
rect 108684 386280 108946 386336
rect 109002 386280 109007 386336
rect 108684 386278 109007 386280
rect 108684 386276 108690 386278
rect 108941 386275 109007 386278
rect 111006 386276 111012 386340
rect 111076 386338 111082 386340
rect 111701 386338 111767 386341
rect 111076 386336 111767 386338
rect 111076 386280 111706 386336
rect 111762 386280 111767 386336
rect 111076 386278 111767 386280
rect 111076 386276 111082 386278
rect 111701 386275 111767 386278
rect 115974 386276 115980 386340
rect 116044 386338 116050 386340
rect 117221 386338 117287 386341
rect 118601 386340 118667 386341
rect 116044 386336 117287 386338
rect 116044 386280 117226 386336
rect 117282 386280 117287 386336
rect 116044 386278 117287 386280
rect 116044 386276 116050 386278
rect 117221 386275 117287 386278
rect 118550 386276 118556 386340
rect 118620 386338 118667 386340
rect 118620 386336 118712 386338
rect 118662 386280 118712 386336
rect 118620 386278 118712 386280
rect 118620 386276 118667 386278
rect 123518 386276 123524 386340
rect 123588 386338 123594 386340
rect 124121 386338 124187 386341
rect 123588 386336 124187 386338
rect 123588 386280 124126 386336
rect 124182 386280 124187 386336
rect 123588 386278 124187 386280
rect 123588 386276 123594 386278
rect 118601 386275 118667 386276
rect 124121 386275 124187 386278
rect 125910 386276 125916 386340
rect 125980 386338 125986 386340
rect 126881 386338 126947 386341
rect 133689 386340 133755 386341
rect 138473 386340 138539 386341
rect 133638 386338 133644 386340
rect 125980 386336 126947 386338
rect 125980 386280 126886 386336
rect 126942 386280 126947 386336
rect 125980 386278 126947 386280
rect 133598 386278 133644 386338
rect 133708 386336 133755 386340
rect 138422 386338 138428 386340
rect 133750 386280 133755 386336
rect 125980 386276 125986 386278
rect 126881 386275 126947 386278
rect 133638 386276 133644 386278
rect 133708 386276 133755 386280
rect 138382 386278 138428 386338
rect 138492 386336 138539 386340
rect 138534 386280 138539 386336
rect 138422 386276 138428 386278
rect 138492 386276 138539 386280
rect 140998 386276 141004 386340
rect 141068 386338 141074 386340
rect 142061 386338 142127 386341
rect 143441 386340 143507 386341
rect 158529 386340 158595 386341
rect 159817 386340 159883 386341
rect 143390 386338 143396 386340
rect 141068 386336 142127 386338
rect 141068 386280 142066 386336
rect 142122 386280 142127 386336
rect 141068 386278 142127 386280
rect 143350 386278 143396 386338
rect 143460 386336 143507 386340
rect 158478 386338 158484 386340
rect 143502 386280 143507 386336
rect 141068 386276 141074 386278
rect 133689 386275 133755 386276
rect 138473 386275 138539 386276
rect 142061 386275 142127 386278
rect 143390 386276 143396 386278
rect 143460 386276 143507 386280
rect 158438 386278 158484 386338
rect 158548 386336 158595 386340
rect 159766 386338 159772 386340
rect 158590 386280 158595 386336
rect 158478 386276 158484 386278
rect 158548 386276 158595 386280
rect 159726 386278 159772 386338
rect 159836 386336 159883 386340
rect 159878 386280 159883 386336
rect 159766 386276 159772 386278
rect 159836 386276 159883 386280
rect 143441 386275 143507 386276
rect 158529 386275 158595 386276
rect 159817 386275 159883 386276
rect 248505 386338 248571 386341
rect 248638 386338 248644 386340
rect 248505 386336 248644 386338
rect 248505 386280 248510 386336
rect 248566 386280 248644 386336
rect 248505 386278 248644 386280
rect 248505 386275 248571 386278
rect 248638 386276 248644 386278
rect 248708 386276 248714 386340
rect 252553 386338 252619 386341
rect 253422 386338 253428 386340
rect 252553 386336 253428 386338
rect 252553 386280 252558 386336
rect 252614 386280 253428 386336
rect 252553 386278 253428 386280
rect 252553 386275 252619 386278
rect 253422 386276 253428 386278
rect 253492 386276 253498 386340
rect 255313 386338 255379 386341
rect 256182 386338 256188 386340
rect 255313 386336 256188 386338
rect 255313 386280 255318 386336
rect 255374 386280 256188 386336
rect 255313 386278 256188 386280
rect 255313 386275 255379 386278
rect 256182 386276 256188 386278
rect 256252 386276 256258 386340
rect 258257 386338 258323 386341
rect 258390 386338 258396 386340
rect 258257 386336 258396 386338
rect 258257 386280 258262 386336
rect 258318 386280 258396 386336
rect 258257 386278 258396 386280
rect 258257 386275 258323 386278
rect 258390 386276 258396 386278
rect 258460 386276 258466 386340
rect 260833 386338 260899 386341
rect 263593 386340 263659 386341
rect 260966 386338 260972 386340
rect 260833 386336 260972 386338
rect 260833 386280 260838 386336
rect 260894 386280 260972 386336
rect 260833 386278 260972 386280
rect 260833 386275 260899 386278
rect 260966 386276 260972 386278
rect 261036 386276 261042 386340
rect 263542 386276 263548 386340
rect 263612 386338 263659 386340
rect 264973 386338 265039 386341
rect 266118 386338 266124 386340
rect 263612 386336 263704 386338
rect 263654 386280 263704 386336
rect 263612 386278 263704 386280
rect 264973 386336 266124 386338
rect 264973 386280 264978 386336
rect 265034 386280 266124 386336
rect 264973 386278 266124 386280
rect 263612 386276 263659 386278
rect 263593 386275 263659 386276
rect 264973 386275 265039 386278
rect 266118 386276 266124 386278
rect 266188 386276 266194 386340
rect 268101 386338 268167 386341
rect 268510 386338 268516 386340
rect 268101 386336 268516 386338
rect 268101 386280 268106 386336
rect 268162 386280 268516 386336
rect 268101 386278 268516 386280
rect 268101 386275 268167 386278
rect 268510 386276 268516 386278
rect 268580 386276 268586 386340
rect 270493 386338 270559 386341
rect 271086 386338 271092 386340
rect 270493 386336 271092 386338
rect 270493 386280 270498 386336
rect 270554 386280 271092 386336
rect 270493 386278 271092 386280
rect 270493 386275 270559 386278
rect 271086 386276 271092 386278
rect 271156 386276 271162 386340
rect 273253 386338 273319 386341
rect 273478 386338 273484 386340
rect 273253 386336 273484 386338
rect 273253 386280 273258 386336
rect 273314 386280 273484 386336
rect 273253 386278 273484 386280
rect 273253 386275 273319 386278
rect 273478 386276 273484 386278
rect 273548 386276 273554 386340
rect 277945 386338 278011 386341
rect 278446 386338 278452 386340
rect 277945 386336 278452 386338
rect 277945 386280 277950 386336
rect 278006 386280 278452 386336
rect 277945 386278 278452 386280
rect 277945 386275 278011 386278
rect 278446 386276 278452 386278
rect 278516 386276 278522 386340
rect 280153 386338 280219 386341
rect 280838 386338 280844 386340
rect 280153 386336 280844 386338
rect 280153 386280 280158 386336
rect 280214 386280 280844 386336
rect 280153 386278 280844 386280
rect 280153 386275 280219 386278
rect 280838 386276 280844 386278
rect 280908 386276 280914 386340
rect 288433 386338 288499 386341
rect 288566 386338 288572 386340
rect 288433 386336 288572 386338
rect 288433 386280 288438 386336
rect 288494 386280 288572 386336
rect 288433 386278 288572 386280
rect 288433 386275 288499 386278
rect 288566 386276 288572 386278
rect 288636 386276 288642 386340
rect 295333 386338 295399 386341
rect 295926 386338 295932 386340
rect 295333 386336 295932 386338
rect 295333 386280 295338 386336
rect 295394 386280 295932 386336
rect 295333 386278 295932 386280
rect 295333 386275 295399 386278
rect 295926 386276 295932 386278
rect 295996 386276 296002 386340
rect 304993 386338 305059 386341
rect 305862 386338 305868 386340
rect 304993 386336 305868 386338
rect 304993 386280 304998 386336
rect 305054 386280 305868 386336
rect 304993 386278 305868 386280
rect 304993 386275 305059 386278
rect 305862 386276 305868 386278
rect 305932 386276 305938 386340
rect 310513 386338 310579 386341
rect 311014 386338 311020 386340
rect 310513 386336 311020 386338
rect 310513 386280 310518 386336
rect 310574 386280 311020 386336
rect 310513 386278 311020 386280
rect 310513 386275 310579 386278
rect 311014 386276 311020 386278
rect 311084 386276 311090 386340
rect 313273 386338 313339 386341
rect 313590 386338 313596 386340
rect 313273 386336 313596 386338
rect 313273 386280 313278 386336
rect 313334 386280 313596 386336
rect 313273 386278 313596 386280
rect 313273 386275 313339 386278
rect 313590 386276 313596 386278
rect 313660 386276 313666 386340
rect 317413 386338 317479 386341
rect 318374 386338 318380 386340
rect 317413 386336 318380 386338
rect 317413 386280 317418 386336
rect 317474 386280 318380 386336
rect 317413 386278 318380 386280
rect 317413 386275 317479 386278
rect 318374 386276 318380 386278
rect 318444 386276 318450 386340
rect 320173 386338 320239 386341
rect 320950 386338 320956 386340
rect 320173 386336 320956 386338
rect 320173 386280 320178 386336
rect 320234 386280 320956 386336
rect 320173 386278 320956 386280
rect 320173 386275 320239 386278
rect 320950 386276 320956 386278
rect 321020 386276 321026 386340
rect 322933 386338 322999 386341
rect 323342 386338 323348 386340
rect 322933 386336 323348 386338
rect 322933 386280 322938 386336
rect 322994 386280 323348 386336
rect 322933 386278 323348 386280
rect 322933 386275 322999 386278
rect 323342 386276 323348 386278
rect 323412 386276 323418 386340
rect 338113 386338 338179 386341
rect 338430 386338 338436 386340
rect 338113 386336 338436 386338
rect 338113 386280 338118 386336
rect 338174 386280 338436 386336
rect 338113 386278 338436 386280
rect 338113 386275 338179 386278
rect 338430 386276 338436 386278
rect 338500 386276 338506 386340
rect 339493 386338 339559 386341
rect 339718 386338 339724 386340
rect 339493 386336 339724 386338
rect 339493 386280 339498 386336
rect 339554 386280 339724 386336
rect 339493 386278 339724 386280
rect 339493 386275 339559 386278
rect 339718 386276 339724 386278
rect 339788 386276 339794 386340
rect 285673 386202 285739 386205
rect 285990 386202 285996 386204
rect 285673 386200 285996 386202
rect 285673 386144 285678 386200
rect 285734 386144 285996 386200
rect 285673 386142 285996 386144
rect 285673 386139 285739 386142
rect 285990 386140 285996 386142
rect 286060 386140 286066 386204
rect 289813 386202 289879 386205
rect 290958 386202 290964 386204
rect 289813 386200 290964 386202
rect 289813 386144 289818 386200
rect 289874 386144 290964 386200
rect 289813 386142 290964 386144
rect 289813 386139 289879 386142
rect 290958 386140 290964 386142
rect 291028 386140 291034 386204
rect 249793 386066 249859 386069
rect 251030 386066 251036 386068
rect 249793 386064 251036 386066
rect 249793 386008 249798 386064
rect 249854 386008 251036 386064
rect 249793 386006 251036 386008
rect 249793 386003 249859 386006
rect 251030 386004 251036 386006
rect 251100 386004 251106 386068
rect 316033 386066 316099 386069
rect 316166 386066 316172 386068
rect 316033 386064 316172 386066
rect 316033 386008 316038 386064
rect 316094 386008 316172 386064
rect 316033 386006 316172 386008
rect 316033 386003 316099 386006
rect 316166 386004 316172 386006
rect 316236 386004 316242 386068
rect 298093 385930 298159 385933
rect 298502 385930 298508 385932
rect 298093 385928 298508 385930
rect 298093 385872 298098 385928
rect 298154 385872 298508 385928
rect 298093 385870 298508 385872
rect 298093 385867 298159 385870
rect 298502 385868 298508 385870
rect 298572 385868 298578 385932
rect 302233 385930 302299 385933
rect 303470 385930 303476 385932
rect 302233 385928 303476 385930
rect 302233 385872 302238 385928
rect 302294 385872 303476 385928
rect 302233 385870 303476 385872
rect 302233 385867 302299 385870
rect 303470 385868 303476 385870
rect 303540 385868 303546 385932
rect 103646 385188 103652 385252
rect 103716 385250 103722 385252
rect 104801 385250 104867 385253
rect 103716 385248 104867 385250
rect 103716 385192 104806 385248
rect 104862 385192 104867 385248
rect 103716 385190 104867 385192
rect 103716 385188 103722 385190
rect 104801 385187 104867 385190
rect 73470 385052 73476 385116
rect 73540 385114 73546 385116
rect 73889 385114 73955 385117
rect 73540 385112 73955 385114
rect 73540 385056 73894 385112
rect 73950 385056 73955 385112
rect 73540 385054 73955 385056
rect 73540 385052 73546 385054
rect 73889 385051 73955 385054
rect 76230 385052 76236 385116
rect 76300 385114 76306 385116
rect 77201 385114 77267 385117
rect 81065 385116 81131 385117
rect 83641 385116 83707 385117
rect 81014 385114 81020 385116
rect 76300 385112 77267 385114
rect 76300 385056 77206 385112
rect 77262 385056 77267 385112
rect 76300 385054 77267 385056
rect 80974 385054 81020 385114
rect 81084 385112 81131 385116
rect 83590 385114 83596 385116
rect 81126 385056 81131 385112
rect 76300 385052 76306 385054
rect 77201 385051 77267 385054
rect 81014 385052 81020 385054
rect 81084 385052 81131 385056
rect 83550 385054 83596 385114
rect 83660 385112 83707 385116
rect 83702 385056 83707 385112
rect 83590 385052 83596 385054
rect 83660 385052 83707 385056
rect 86166 385052 86172 385116
rect 86236 385114 86242 385116
rect 86493 385114 86559 385117
rect 86236 385112 86559 385114
rect 86236 385056 86498 385112
rect 86554 385056 86559 385112
rect 86236 385054 86559 385056
rect 86236 385052 86242 385054
rect 81065 385051 81131 385052
rect 83641 385051 83707 385052
rect 86493 385051 86559 385054
rect 91134 385052 91140 385116
rect 91204 385114 91210 385116
rect 92105 385114 92171 385117
rect 91204 385112 92171 385114
rect 91204 385056 92110 385112
rect 92166 385056 92171 385112
rect 91204 385054 92171 385056
rect 91204 385052 91210 385054
rect 92105 385051 92171 385054
rect 113582 385052 113588 385116
rect 113652 385114 113658 385116
rect 114461 385114 114527 385117
rect 113652 385112 114527 385114
rect 113652 385056 114466 385112
rect 114522 385056 114527 385112
rect 113652 385054 114527 385056
rect 113652 385052 113658 385054
rect 114461 385051 114527 385054
rect 121126 385052 121132 385116
rect 121196 385114 121202 385116
rect 121361 385114 121427 385117
rect 121196 385112 121427 385114
rect 121196 385056 121366 385112
rect 121422 385056 121427 385112
rect 121196 385054 121427 385056
rect 121196 385052 121202 385054
rect 121361 385051 121427 385054
rect 128486 385052 128492 385116
rect 128556 385114 128562 385116
rect 128629 385114 128695 385117
rect 128556 385112 128695 385114
rect 128556 385056 128634 385112
rect 128690 385056 128695 385112
rect 128556 385054 128695 385056
rect 128556 385052 128562 385054
rect 128629 385051 128695 385054
rect 131021 385116 131087 385117
rect 136081 385116 136147 385117
rect 146201 385116 146267 385117
rect 131021 385112 131068 385116
rect 131132 385114 131138 385116
rect 136030 385114 136036 385116
rect 131021 385056 131026 385112
rect 131021 385052 131068 385056
rect 131132 385054 131178 385114
rect 135990 385054 136036 385114
rect 136100 385112 136147 385116
rect 146150 385114 146156 385116
rect 136142 385056 136147 385112
rect 131132 385052 131138 385054
rect 136030 385052 136036 385054
rect 136100 385052 136147 385056
rect 146110 385054 146156 385114
rect 146220 385112 146267 385116
rect 276013 385116 276079 385117
rect 276013 385114 276060 385116
rect 146262 385056 146267 385112
rect 146150 385052 146156 385054
rect 146220 385052 146267 385056
rect 275968 385112 276060 385114
rect 275968 385056 276018 385112
rect 275968 385054 276060 385056
rect 131021 385051 131087 385052
rect 136081 385051 136147 385052
rect 146201 385051 146267 385052
rect 276013 385052 276060 385054
rect 276124 385052 276130 385116
rect 282913 385114 282979 385117
rect 283598 385114 283604 385116
rect 282913 385112 283604 385114
rect 282913 385056 282918 385112
rect 282974 385056 283604 385112
rect 282913 385054 283604 385056
rect 276013 385051 276079 385052
rect 282913 385051 282979 385054
rect 283598 385052 283604 385054
rect 283668 385052 283674 385116
rect 292573 385114 292639 385117
rect 293534 385114 293540 385116
rect 292573 385112 293540 385114
rect 292573 385056 292578 385112
rect 292634 385056 293540 385112
rect 292573 385054 293540 385056
rect 292573 385051 292639 385054
rect 293534 385052 293540 385054
rect 293604 385052 293610 385116
rect 300853 385114 300919 385117
rect 301078 385114 301084 385116
rect 300853 385112 301084 385114
rect 300853 385056 300858 385112
rect 300914 385056 301084 385112
rect 300853 385054 301084 385056
rect 300853 385051 300919 385054
rect 301078 385052 301084 385054
rect 301148 385052 301154 385116
rect 307753 385114 307819 385117
rect 308438 385114 308444 385116
rect 307753 385112 308444 385114
rect 307753 385056 307758 385112
rect 307814 385056 308444 385112
rect 307753 385054 308444 385056
rect 307753 385051 307819 385054
rect 308438 385052 308444 385054
rect 308508 385052 308514 385116
rect 325877 385114 325943 385117
rect 350993 385116 351059 385117
rect 326102 385114 326108 385116
rect 325877 385112 326108 385114
rect 325877 385056 325882 385112
rect 325938 385056 326108 385112
rect 325877 385054 326108 385056
rect 325877 385051 325943 385054
rect 326102 385052 326108 385054
rect 326172 385052 326178 385116
rect 350942 385114 350948 385116
rect 350902 385054 350948 385114
rect 351012 385112 351059 385116
rect 351054 385056 351059 385112
rect 350942 385052 350948 385054
rect 351012 385052 351059 385056
rect 350993 385051 351059 385052
rect -960 384284 480 384524
rect 170857 384164 170923 384165
rect 170806 384162 170812 384164
rect 170766 384102 170812 384162
rect 170876 384160 170923 384164
rect 170918 384104 170923 384160
rect 170806 384100 170812 384102
rect 170876 384100 170923 384104
rect 170857 384099 170923 384100
rect 359273 379402 359339 379405
rect 356562 379400 359339 379402
rect 356562 379344 359278 379400
rect 359334 379344 359339 379400
rect 356562 379342 359339 379344
rect 178677 379266 178743 379269
rect 177070 379264 178743 379266
rect 177070 379220 178682 379264
rect 176548 379208 178682 379220
rect 178738 379208 178743 379264
rect 176548 379206 178743 379208
rect 176548 379160 177130 379206
rect 178677 379203 178743 379206
rect 356562 379190 356622 379342
rect 359273 379339 359339 379342
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect 38285 336834 38351 336837
rect 39990 336834 40050 336894
rect 219390 336864 220064 336924
rect 38285 336832 40050 336834
rect 38285 336776 38290 336832
rect 38346 336776 40050 336832
rect 38285 336774 40050 336776
rect 216673 336834 216739 336837
rect 219390 336834 219450 336864
rect 216673 336832 219450 336834
rect 216673 336776 216678 336832
rect 216734 336776 219450 336832
rect 216673 336774 219450 336776
rect 38285 336771 38351 336774
rect 216673 336771 216739 336774
rect 38745 335610 38811 335613
rect 39990 335610 40050 335942
rect 219390 335912 220064 335972
rect 217317 335882 217383 335885
rect 219390 335882 219450 335912
rect 217317 335880 219450 335882
rect 217317 335824 217322 335880
rect 217378 335824 219450 335880
rect 217317 335822 219450 335824
rect 217317 335819 217383 335822
rect 38745 335608 40050 335610
rect 38745 335552 38750 335608
rect 38806 335552 40050 335608
rect 38745 335550 40050 335552
rect 38745 335547 38811 335550
rect 38377 333162 38443 333165
rect 39990 333162 40050 333766
rect 219390 333736 220064 333796
rect 217961 333706 218027 333709
rect 219390 333706 219450 333736
rect 217961 333704 219450 333706
rect 217961 333648 217966 333704
rect 218022 333648 219450 333704
rect 217961 333646 219450 333648
rect 217961 333643 218027 333646
rect 38377 333160 40050 333162
rect 38377 333104 38382 333160
rect 38438 333104 40050 333160
rect 38377 333102 40050 333104
rect 38377 333099 38443 333102
rect 38561 332618 38627 332621
rect 39990 332618 40050 332814
rect 219390 332784 220064 332844
rect 217542 332692 217548 332756
rect 217612 332754 217618 332756
rect 219390 332754 219450 332784
rect 217612 332694 219450 332754
rect 217612 332692 217618 332694
rect 38561 332616 40050 332618
rect 38561 332560 38566 332616
rect 38622 332560 40050 332616
rect 38561 332558 40050 332560
rect 38561 332555 38627 332558
rect -960 332196 480 332436
rect 39021 330442 39087 330445
rect 39990 330442 40050 331046
rect 219390 331016 220064 331076
rect 217358 330924 217364 330988
rect 217428 330986 217434 330988
rect 219390 330986 219450 331016
rect 217428 330926 219450 330986
rect 217428 330924 217434 330926
rect 39021 330440 40050 330442
rect 39021 330384 39026 330440
rect 39082 330384 40050 330440
rect 39021 330382 40050 330384
rect 39021 330379 39087 330382
rect 38837 329898 38903 329901
rect 39990 329898 40050 329958
rect 219390 329928 220064 329988
rect 38837 329896 40050 329898
rect 38837 329840 38842 329896
rect 38898 329840 40050 329896
rect 38837 329838 40050 329840
rect 217501 329898 217567 329901
rect 219390 329898 219450 329928
rect 217501 329896 219450 329898
rect 217501 329840 217506 329896
rect 217562 329840 219450 329896
rect 217501 329838 219450 329840
rect 38837 329835 38903 329838
rect 217501 329835 217567 329838
rect 38653 327586 38719 327589
rect 39990 327586 40050 328190
rect 219390 328160 220064 328220
rect 217174 328068 217180 328132
rect 217244 328130 217250 328132
rect 219390 328130 219450 328160
rect 217244 328070 219450 328130
rect 217244 328068 217250 328070
rect 38653 327584 40050 327586
rect 38653 327528 38658 327584
rect 38714 327528 40050 327584
rect 38653 327526 40050 327528
rect 38653 327523 38719 327526
rect 583520 325124 584960 325364
rect 359181 319970 359247 319973
rect 356562 319968 359247 319970
rect 356562 319912 359186 319968
rect 359242 319912 359247 319968
rect 356562 319910 359247 319912
rect 178677 319426 178743 319429
rect 177070 319424 178743 319426
rect 177070 319380 178682 319424
rect -960 319140 480 319380
rect 176548 319368 178682 319380
rect 178738 319368 178743 319424
rect 176548 319366 178743 319368
rect 176548 319320 177130 319366
rect 178677 319363 178743 319366
rect 356562 319350 356622 319910
rect 359181 319907 359247 319910
rect 359089 318338 359155 318341
rect 356562 318336 359155 318338
rect 356562 318280 359094 318336
rect 359150 318280 359155 318336
rect 356562 318278 359155 318280
rect 178953 317794 179019 317797
rect 177070 317792 179019 317794
rect 177070 317748 178958 317792
rect 176548 317736 178958 317748
rect 179014 317736 179019 317792
rect 176548 317734 179019 317736
rect 176548 317688 177130 317734
rect 178953 317731 179019 317734
rect 356562 317718 356622 318278
rect 359089 318275 359155 318278
rect 358997 316978 359063 316981
rect 356562 316976 359063 316978
rect 356562 316920 359002 316976
rect 359058 316920 359063 316976
rect 356562 316918 359063 316920
rect 178953 316434 179019 316437
rect 177070 316432 179019 316434
rect 177070 316388 178958 316432
rect 176548 316376 178958 316388
rect 179014 316376 179019 316432
rect 176548 316374 179019 316376
rect 176548 316328 177130 316374
rect 178953 316371 179019 316374
rect 356562 316358 356622 316918
rect 358997 316915 359063 316918
rect 358905 315482 358971 315485
rect 356562 315480 358971 315482
rect 356562 315424 358910 315480
rect 358966 315424 358971 315480
rect 356562 315422 358971 315424
rect 178585 314938 178651 314941
rect 177070 314936 178651 314938
rect 177070 314892 178590 314936
rect 176548 314880 178590 314892
rect 178646 314880 178651 314936
rect 176548 314878 178651 314880
rect 176548 314832 177130 314878
rect 178585 314875 178651 314878
rect 356562 314862 356622 315422
rect 358905 315419 358971 315422
rect 358813 314258 358879 314261
rect 356562 314256 358879 314258
rect 356562 314200 358818 314256
rect 358874 314200 358879 314256
rect 356562 314198 358879 314200
rect 178677 313714 178743 313717
rect 177070 313712 178743 313714
rect 177070 313668 178682 313712
rect 176548 313656 178682 313668
rect 178738 313656 178743 313712
rect 176548 313654 178743 313656
rect 176548 313608 177130 313654
rect 178677 313651 178743 313654
rect 356562 313638 356622 314198
rect 358813 314195 358879 314198
rect 583520 311932 584960 312172
rect 38469 309362 38535 309365
rect 39990 309362 40050 309966
rect 219390 309936 220064 309996
rect 216673 309906 216739 309909
rect 219390 309906 219450 309936
rect 216673 309904 219450 309906
rect 216673 309848 216678 309904
rect 216734 309848 219450 309904
rect 216673 309846 219450 309848
rect 216673 309843 216739 309846
rect 38469 309360 40050 309362
rect 38469 309304 38474 309360
rect 38530 309304 40050 309360
rect 38469 309302 40050 309304
rect 38469 309299 38535 309302
rect 39113 308410 39179 308413
rect 216765 308410 216831 308413
rect 217869 308410 217935 308413
rect 39113 308408 40050 308410
rect 39113 308352 39118 308408
rect 39174 308352 40050 308408
rect 39113 308350 40050 308352
rect 39113 308347 39179 308350
rect 39990 308334 40050 308350
rect 216765 308408 219450 308410
rect 216765 308352 216770 308408
rect 216826 308352 217874 308408
rect 217930 308364 219450 308408
rect 217930 308352 220064 308364
rect 216765 308350 220064 308352
rect 216765 308347 216831 308350
rect 217869 308347 217935 308350
rect 219390 308304 220064 308350
rect 38929 307866 38995 307869
rect 39990 307866 40050 308062
rect 219390 308032 220064 308092
rect 217869 308002 217935 308005
rect 219390 308002 219450 308032
rect 217869 308000 219450 308002
rect 217869 307944 217874 308000
rect 217930 307944 219450 308000
rect 217869 307942 219450 307944
rect 217869 307939 217935 307942
rect 38929 307864 40050 307866
rect 38929 307808 38934 307864
rect 38990 307808 40050 307864
rect 38929 307806 40050 307808
rect 38929 307803 38995 307806
rect -960 306084 480 306324
rect 163221 299572 163287 299573
rect 163405 299572 163471 299573
rect 163216 299570 163222 299572
rect 163130 299510 163222 299570
rect 163216 299508 163222 299510
rect 163286 299508 163292 299572
rect 163352 299508 163358 299572
rect 163422 299570 163471 299572
rect 163422 299568 163514 299570
rect 163466 299512 163514 299568
rect 163422 299510 163514 299512
rect 163422 299508 163471 299510
rect 163221 299507 163287 299508
rect 163405 299507 163471 299508
rect 583520 298604 584960 298844
rect 55990 298148 55996 298212
rect 56060 298148 56066 298212
rect 59670 298148 59676 298212
rect 59740 298148 59746 298212
rect 63166 298148 63172 298212
rect 63236 298148 63242 298212
rect 73654 298148 73660 298212
rect 73724 298148 73730 298212
rect 85246 298148 85252 298212
rect 85316 298148 85322 298212
rect 92238 298148 92244 298212
rect 92308 298148 92314 298212
rect 95734 298148 95740 298212
rect 95804 298148 95810 298212
rect 113398 298148 113404 298212
rect 113468 298148 113474 298212
rect 120942 298148 120948 298212
rect 121012 298148 121018 298212
rect 145966 298148 145972 298212
rect 146036 298148 146042 298212
rect 258022 298148 258028 298212
rect 258092 298148 258098 298212
rect 261702 298148 261708 298212
rect 261772 298148 261778 298212
rect 265198 298148 265204 298212
rect 265268 298148 265274 298212
rect 272190 298148 272196 298212
rect 272260 298148 272266 298212
rect 275686 298148 275692 298212
rect 275756 298148 275762 298212
rect 276054 298148 276060 298212
rect 276124 298148 276130 298212
rect 283414 298148 283420 298212
rect 283484 298148 283490 298212
rect 300894 298148 300900 298212
rect 300964 298148 300970 298212
rect 315798 298148 315804 298212
rect 315868 298148 315874 298212
rect 325918 298148 325924 298212
rect 325988 298148 325994 298212
rect 55998 298074 56058 298148
rect 56501 298074 56567 298077
rect 55998 298072 56567 298074
rect 55998 298016 56506 298072
rect 56562 298016 56567 298072
rect 55998 298014 56567 298016
rect 56501 298011 56567 298014
rect 57094 298012 57100 298076
rect 57164 298074 57170 298076
rect 57881 298074 57947 298077
rect 57164 298072 57947 298074
rect 57164 298016 57886 298072
rect 57942 298016 57947 298072
rect 57164 298014 57947 298016
rect 57164 298012 57170 298014
rect 57881 298011 57947 298014
rect 58198 298012 58204 298076
rect 58268 298074 58274 298076
rect 59261 298074 59327 298077
rect 58268 298072 59327 298074
rect 58268 298016 59266 298072
rect 59322 298016 59327 298072
rect 58268 298014 59327 298016
rect 58268 298012 58274 298014
rect 59261 298011 59327 298014
rect 59678 297938 59738 298148
rect 60641 298076 60707 298077
rect 60590 298074 60596 298076
rect 60550 298014 60596 298074
rect 60660 298072 60707 298076
rect 60702 298016 60707 298072
rect 60590 298012 60596 298014
rect 60660 298012 60707 298016
rect 61878 298012 61884 298076
rect 61948 298074 61954 298076
rect 62021 298074 62087 298077
rect 61948 298072 62087 298074
rect 61948 298016 62026 298072
rect 62082 298016 62087 298072
rect 61948 298014 62087 298016
rect 63174 298074 63234 298148
rect 63401 298074 63467 298077
rect 63174 298072 63467 298074
rect 63174 298016 63406 298072
rect 63462 298016 63467 298072
rect 63174 298014 63467 298016
rect 61948 298012 61954 298014
rect 60641 298011 60707 298012
rect 62021 298011 62087 298014
rect 63401 298011 63467 298014
rect 64270 298012 64276 298076
rect 64340 298074 64346 298076
rect 64781 298074 64847 298077
rect 64340 298072 64847 298074
rect 64340 298016 64786 298072
rect 64842 298016 64847 298072
rect 64340 298014 64847 298016
rect 64340 298012 64346 298014
rect 64781 298011 64847 298014
rect 65374 298012 65380 298076
rect 65444 298074 65450 298076
rect 66161 298074 66227 298077
rect 65444 298072 66227 298074
rect 65444 298016 66166 298072
rect 66222 298016 66227 298072
rect 65444 298014 66227 298016
rect 65444 298012 65450 298014
rect 66161 298011 66227 298014
rect 66478 298012 66484 298076
rect 66548 298074 66554 298076
rect 67541 298074 67607 298077
rect 66548 298072 67607 298074
rect 66548 298016 67546 298072
rect 67602 298016 67607 298072
rect 66548 298014 67607 298016
rect 66548 298012 66554 298014
rect 67541 298011 67607 298014
rect 68318 298012 68324 298076
rect 68388 298074 68394 298076
rect 68737 298074 68803 298077
rect 68388 298072 68803 298074
rect 68388 298016 68742 298072
rect 68798 298016 68803 298072
rect 68388 298014 68803 298016
rect 68388 298012 68394 298014
rect 68737 298011 68803 298014
rect 70158 298012 70164 298076
rect 70228 298074 70234 298076
rect 70301 298074 70367 298077
rect 70228 298072 70367 298074
rect 70228 298016 70306 298072
rect 70362 298016 70367 298072
rect 70228 298014 70367 298016
rect 70228 298012 70234 298014
rect 70301 298011 70367 298014
rect 71262 298012 71268 298076
rect 71332 298074 71338 298076
rect 71681 298074 71747 298077
rect 71332 298072 71747 298074
rect 71332 298016 71686 298072
rect 71742 298016 71747 298072
rect 71332 298014 71747 298016
rect 71332 298012 71338 298014
rect 71681 298011 71747 298014
rect 72366 298012 72372 298076
rect 72436 298074 72442 298076
rect 73061 298074 73127 298077
rect 72436 298072 73127 298074
rect 72436 298016 73066 298072
rect 73122 298016 73127 298072
rect 72436 298014 73127 298016
rect 73662 298074 73722 298148
rect 74441 298074 74507 298077
rect 73662 298072 74507 298074
rect 73662 298016 74446 298072
rect 74502 298016 74507 298072
rect 73662 298014 74507 298016
rect 72436 298012 72442 298014
rect 73061 298011 73127 298014
rect 74441 298011 74507 298014
rect 74574 298012 74580 298076
rect 74644 298074 74650 298076
rect 75821 298074 75887 298077
rect 74644 298072 75887 298074
rect 74644 298016 75826 298072
rect 75882 298016 75887 298072
rect 74644 298014 75887 298016
rect 74644 298012 74650 298014
rect 75821 298011 75887 298014
rect 76046 298012 76052 298076
rect 76116 298074 76122 298076
rect 77017 298074 77083 298077
rect 78489 298076 78555 298077
rect 78438 298074 78444 298076
rect 76116 298072 77083 298074
rect 76116 298016 77022 298072
rect 77078 298016 77083 298072
rect 76116 298014 77083 298016
rect 78398 298014 78444 298074
rect 78508 298072 78555 298076
rect 78550 298016 78555 298072
rect 76116 298012 76122 298014
rect 77017 298011 77083 298014
rect 78438 298012 78444 298014
rect 78508 298012 78555 298016
rect 79542 298012 79548 298076
rect 79612 298074 79618 298076
rect 79961 298074 80027 298077
rect 80697 298076 80763 298077
rect 80646 298074 80652 298076
rect 79612 298072 80027 298074
rect 79612 298016 79966 298072
rect 80022 298016 80027 298072
rect 79612 298014 80027 298016
rect 80606 298014 80652 298074
rect 80716 298072 80763 298076
rect 80758 298016 80763 298072
rect 79612 298012 79618 298014
rect 78489 298011 78555 298012
rect 79961 298011 80027 298014
rect 80646 298012 80652 298014
rect 80716 298012 80763 298016
rect 81014 298012 81020 298076
rect 81084 298074 81090 298076
rect 81249 298074 81315 298077
rect 81084 298072 81315 298074
rect 81084 298016 81254 298072
rect 81310 298016 81315 298072
rect 81084 298014 81315 298016
rect 81084 298012 81090 298014
rect 80697 298011 80763 298012
rect 81249 298011 81315 298014
rect 81934 298012 81940 298076
rect 82004 298074 82010 298076
rect 82721 298074 82787 298077
rect 82004 298072 82787 298074
rect 82004 298016 82726 298072
rect 82782 298016 82787 298072
rect 82004 298014 82787 298016
rect 82004 298012 82010 298014
rect 82721 298011 82787 298014
rect 82854 298012 82860 298076
rect 82924 298074 82930 298076
rect 83365 298074 83431 298077
rect 84009 298076 84075 298077
rect 83958 298074 83964 298076
rect 82924 298072 83431 298074
rect 82924 298016 83370 298072
rect 83426 298016 83431 298072
rect 82924 298014 83431 298016
rect 83918 298014 83964 298074
rect 84028 298072 84075 298076
rect 84070 298016 84075 298072
rect 82924 298012 82930 298014
rect 83365 298011 83431 298014
rect 83958 298012 83964 298014
rect 84028 298012 84075 298016
rect 85254 298074 85314 298148
rect 85481 298074 85547 298077
rect 85254 298072 85547 298074
rect 85254 298016 85486 298072
rect 85542 298016 85547 298072
rect 85254 298014 85547 298016
rect 84009 298011 84075 298012
rect 85481 298011 85547 298014
rect 85982 298012 85988 298076
rect 86052 298074 86058 298076
rect 86217 298074 86283 298077
rect 86052 298072 86283 298074
rect 86052 298016 86222 298072
rect 86278 298016 86283 298072
rect 86052 298014 86283 298016
rect 86052 298012 86058 298014
rect 86217 298011 86283 298014
rect 86350 298012 86356 298076
rect 86420 298074 86426 298076
rect 86769 298074 86835 298077
rect 86420 298072 86835 298074
rect 86420 298016 86774 298072
rect 86830 298016 86835 298072
rect 86420 298014 86835 298016
rect 86420 298012 86426 298014
rect 86769 298011 86835 298014
rect 88149 298076 88215 298077
rect 88149 298072 88196 298076
rect 88260 298074 88266 298076
rect 88149 298016 88154 298072
rect 88149 298012 88196 298016
rect 88260 298014 88306 298074
rect 88260 298012 88266 298014
rect 88742 298012 88748 298076
rect 88812 298074 88818 298076
rect 89621 298074 89687 298077
rect 91001 298076 91067 298077
rect 90950 298074 90956 298076
rect 88812 298072 89687 298074
rect 88812 298016 89626 298072
rect 89682 298016 89687 298072
rect 88812 298014 89687 298016
rect 90910 298014 90956 298074
rect 91020 298072 91067 298076
rect 91062 298016 91067 298072
rect 88812 298012 88818 298014
rect 88149 298011 88215 298012
rect 89621 298011 89687 298014
rect 90950 298012 90956 298014
rect 91020 298012 91067 298016
rect 92246 298074 92306 298148
rect 92381 298074 92447 298077
rect 92246 298072 92447 298074
rect 92246 298016 92386 298072
rect 92442 298016 92447 298072
rect 92246 298014 92447 298016
rect 91001 298011 91067 298012
rect 92381 298011 92447 298014
rect 93526 298012 93532 298076
rect 93596 298074 93602 298076
rect 93761 298074 93827 298077
rect 93596 298072 93827 298074
rect 93596 298016 93766 298072
rect 93822 298016 93827 298072
rect 93596 298014 93827 298016
rect 93596 298012 93602 298014
rect 93761 298011 93827 298014
rect 94446 298012 94452 298076
rect 94516 298074 94522 298076
rect 95141 298074 95207 298077
rect 94516 298072 95207 298074
rect 94516 298016 95146 298072
rect 95202 298016 95207 298072
rect 94516 298014 95207 298016
rect 94516 298012 94522 298014
rect 95141 298011 95207 298014
rect 60549 297938 60615 297941
rect 59678 297936 60615 297938
rect 59678 297880 60554 297936
rect 60610 297880 60615 297936
rect 59678 297878 60615 297880
rect 60549 297875 60615 297878
rect 68686 297876 68692 297940
rect 68756 297938 68762 297940
rect 68829 297938 68895 297941
rect 68756 297936 68895 297938
rect 68756 297880 68834 297936
rect 68890 297880 68895 297936
rect 68756 297878 68895 297880
rect 68756 297876 68762 297878
rect 68829 297875 68895 297878
rect 73470 297876 73476 297940
rect 73540 297938 73546 297940
rect 74349 297938 74415 297941
rect 73540 297936 74415 297938
rect 73540 297880 74354 297936
rect 74410 297880 74415 297936
rect 73540 297878 74415 297880
rect 73540 297876 73546 297878
rect 74349 297875 74415 297878
rect 75862 297876 75868 297940
rect 75932 297938 75938 297940
rect 77109 297938 77175 297941
rect 75932 297936 77175 297938
rect 75932 297880 77114 297936
rect 77170 297880 77175 297936
rect 75932 297878 77175 297880
rect 75932 297876 75938 297878
rect 77109 297875 77175 297878
rect 78254 297876 78260 297940
rect 78324 297938 78330 297940
rect 78581 297938 78647 297941
rect 78324 297936 78647 297938
rect 78324 297880 78586 297936
rect 78642 297880 78647 297936
rect 78324 297878 78647 297880
rect 78324 297876 78330 297878
rect 78581 297875 78647 297878
rect 87638 297876 87644 297940
rect 87708 297938 87714 297940
rect 88241 297938 88307 297941
rect 87708 297936 88307 297938
rect 87708 297880 88246 297936
rect 88302 297880 88307 297936
rect 87708 297878 88307 297880
rect 87708 297876 87714 297878
rect 88241 297875 88307 297878
rect 89846 297876 89852 297940
rect 89916 297938 89922 297940
rect 90909 297938 90975 297941
rect 89916 297936 90975 297938
rect 89916 297880 90914 297936
rect 90970 297880 90975 297936
rect 89916 297878 90975 297880
rect 89916 297876 89922 297878
rect 90909 297875 90975 297878
rect 91134 297876 91140 297940
rect 91204 297938 91210 297940
rect 92289 297938 92355 297941
rect 91204 297936 92355 297938
rect 91204 297880 92294 297936
rect 92350 297880 92355 297936
rect 91204 297878 92355 297880
rect 91204 297876 91210 297878
rect 92289 297875 92355 297878
rect 93342 297876 93348 297940
rect 93412 297938 93418 297940
rect 93669 297938 93735 297941
rect 93412 297936 93735 297938
rect 93412 297880 93674 297936
rect 93730 297880 93735 297936
rect 93412 297878 93735 297880
rect 95742 297938 95802 298148
rect 96286 298012 96292 298076
rect 96356 298074 96362 298076
rect 96429 298074 96495 298077
rect 96356 298072 96495 298074
rect 96356 298016 96434 298072
rect 96490 298016 96495 298072
rect 96356 298014 96495 298016
rect 96356 298012 96362 298014
rect 96429 298011 96495 298014
rect 97022 298012 97028 298076
rect 97092 298074 97098 298076
rect 97901 298074 97967 298077
rect 97092 298072 97967 298074
rect 97092 298016 97906 298072
rect 97962 298016 97967 298072
rect 97092 298014 97967 298016
rect 97092 298012 97098 298014
rect 97901 298011 97967 298014
rect 99046 298012 99052 298076
rect 99116 298074 99122 298076
rect 99189 298074 99255 298077
rect 99116 298072 99255 298074
rect 99116 298016 99194 298072
rect 99250 298016 99255 298072
rect 99116 298014 99255 298016
rect 99116 298012 99122 298014
rect 99189 298011 99255 298014
rect 100886 298012 100892 298076
rect 100956 298074 100962 298076
rect 102041 298074 102107 298077
rect 100956 298072 102107 298074
rect 100956 298016 102046 298072
rect 102102 298016 102107 298072
rect 100956 298014 102107 298016
rect 100956 298012 100962 298014
rect 102041 298011 102107 298014
rect 106038 298012 106044 298076
rect 106108 298074 106114 298076
rect 106181 298074 106247 298077
rect 106108 298072 106247 298074
rect 106108 298016 106186 298072
rect 106242 298016 106247 298072
rect 106108 298014 106247 298016
rect 106108 298012 106114 298014
rect 106181 298011 106247 298014
rect 108246 298012 108252 298076
rect 108316 298074 108322 298076
rect 108481 298074 108547 298077
rect 108316 298072 108547 298074
rect 108316 298016 108486 298072
rect 108542 298016 108547 298072
rect 108316 298014 108547 298016
rect 108316 298012 108322 298014
rect 108481 298011 108547 298014
rect 111006 298012 111012 298076
rect 111076 298074 111082 298076
rect 111701 298074 111767 298077
rect 111076 298072 111767 298074
rect 111076 298016 111706 298072
rect 111762 298016 111767 298072
rect 111076 298014 111767 298016
rect 113406 298074 113466 298148
rect 114461 298074 114527 298077
rect 113406 298072 114527 298074
rect 113406 298016 114466 298072
rect 114522 298016 114527 298072
rect 113406 298014 114527 298016
rect 111076 298012 111082 298014
rect 111701 298011 111767 298014
rect 114461 298011 114527 298014
rect 115933 298076 115999 298077
rect 115933 298072 115980 298076
rect 116044 298074 116050 298076
rect 117405 298074 117471 298077
rect 118366 298074 118372 298076
rect 115933 298016 115938 298072
rect 115933 298012 115980 298016
rect 116044 298014 116090 298074
rect 117405 298072 118372 298074
rect 117405 298016 117410 298072
rect 117466 298016 118372 298072
rect 117405 298014 118372 298016
rect 116044 298012 116050 298014
rect 115933 298011 115999 298012
rect 117405 298011 117471 298014
rect 118366 298012 118372 298014
rect 118436 298012 118442 298076
rect 120950 298074 121010 298148
rect 121361 298074 121427 298077
rect 120950 298072 121427 298074
rect 120950 298016 121366 298072
rect 121422 298016 121427 298072
rect 120950 298014 121427 298016
rect 121361 298011 121427 298014
rect 123518 298012 123524 298076
rect 123588 298074 123594 298076
rect 124121 298074 124187 298077
rect 123588 298072 124187 298074
rect 123588 298016 124126 298072
rect 124182 298016 124187 298072
rect 123588 298014 124187 298016
rect 123588 298012 123594 298014
rect 124121 298011 124187 298014
rect 125869 298076 125935 298077
rect 125869 298072 125916 298076
rect 125980 298074 125986 298076
rect 125869 298016 125874 298072
rect 125869 298012 125916 298016
rect 125980 298014 126026 298074
rect 125980 298012 125986 298014
rect 128670 298012 128676 298076
rect 128740 298074 128746 298076
rect 129641 298074 129707 298077
rect 128740 298072 129707 298074
rect 128740 298016 129646 298072
rect 129702 298016 129707 298072
rect 128740 298014 129707 298016
rect 128740 298012 128746 298014
rect 125869 298011 125935 298012
rect 129641 298011 129707 298014
rect 133454 298012 133460 298076
rect 133524 298074 133530 298076
rect 133781 298074 133847 298077
rect 136081 298076 136147 298077
rect 136030 298074 136036 298076
rect 133524 298072 133847 298074
rect 133524 298016 133786 298072
rect 133842 298016 133847 298072
rect 133524 298014 133847 298016
rect 135990 298014 136036 298074
rect 136100 298072 136147 298076
rect 136142 298016 136147 298072
rect 133524 298012 133530 298014
rect 133781 298011 133847 298014
rect 136030 298012 136036 298014
rect 136100 298012 136147 298016
rect 138422 298012 138428 298076
rect 138492 298074 138498 298076
rect 139301 298074 139367 298077
rect 141049 298076 141115 298077
rect 140998 298074 141004 298076
rect 138492 298072 139367 298074
rect 138492 298016 139306 298072
rect 139362 298016 139367 298072
rect 138492 298014 139367 298016
rect 140958 298014 141004 298074
rect 141068 298072 141115 298076
rect 141110 298016 141115 298072
rect 138492 298012 138498 298014
rect 136081 298011 136147 298012
rect 139301 298011 139367 298014
rect 140998 298012 141004 298014
rect 141068 298012 141115 298016
rect 145974 298074 146034 298148
rect 146201 298074 146267 298077
rect 145974 298072 146267 298074
rect 145974 298016 146206 298072
rect 146262 298016 146267 298072
rect 145974 298014 146267 298016
rect 141049 298011 141115 298012
rect 146201 298011 146267 298014
rect 235993 298074 236059 298077
rect 238109 298076 238175 298077
rect 237046 298074 237052 298076
rect 235993 298072 237052 298074
rect 235993 298016 235998 298072
rect 236054 298016 237052 298072
rect 235993 298014 237052 298016
rect 235993 298011 236059 298014
rect 237046 298012 237052 298014
rect 237116 298012 237122 298076
rect 238109 298072 238156 298076
rect 238220 298074 238226 298076
rect 238109 298016 238114 298072
rect 238109 298012 238156 298016
rect 238220 298014 238266 298074
rect 238220 298012 238226 298014
rect 241830 298012 241836 298076
rect 241900 298074 241906 298076
rect 242801 298074 242867 298077
rect 241900 298072 242867 298074
rect 241900 298016 242806 298072
rect 242862 298016 242867 298072
rect 241900 298014 242867 298016
rect 241900 298012 241906 298014
rect 238109 298011 238175 298012
rect 242801 298011 242867 298014
rect 247033 298074 247099 298077
rect 247718 298074 247724 298076
rect 247033 298072 247724 298074
rect 247033 298016 247038 298072
rect 247094 298016 247724 298072
rect 247033 298014 247724 298016
rect 247033 298011 247099 298014
rect 247718 298012 247724 298014
rect 247788 298012 247794 298076
rect 248413 298074 248479 298077
rect 248638 298074 248644 298076
rect 248413 298072 248644 298074
rect 248413 298016 248418 298072
rect 248474 298016 248644 298072
rect 248413 298014 248644 298016
rect 248413 298011 248479 298014
rect 248638 298012 248644 298014
rect 248708 298012 248714 298076
rect 249793 298074 249859 298077
rect 250110 298074 250116 298076
rect 249793 298072 250116 298074
rect 249793 298016 249798 298072
rect 249854 298016 250116 298072
rect 249793 298014 250116 298016
rect 249793 298011 249859 298014
rect 250110 298012 250116 298014
rect 250180 298012 250186 298076
rect 250846 298012 250852 298076
rect 250916 298074 250922 298076
rect 251081 298074 251147 298077
rect 250916 298072 251147 298074
rect 250916 298016 251086 298072
rect 251142 298016 251147 298072
rect 250916 298014 251147 298016
rect 250916 298012 250922 298014
rect 251081 298011 251147 298014
rect 251214 298012 251220 298076
rect 251284 298074 251290 298076
rect 251357 298074 251423 298077
rect 251284 298072 251423 298074
rect 251284 298016 251362 298072
rect 251418 298016 251423 298072
rect 251284 298014 251423 298016
rect 251284 298012 251290 298014
rect 251357 298011 251423 298014
rect 251541 298074 251607 298077
rect 252318 298074 252324 298076
rect 251541 298072 252324 298074
rect 251541 298016 251546 298072
rect 251602 298016 252324 298072
rect 251541 298014 252324 298016
rect 251541 298011 251607 298014
rect 252318 298012 252324 298014
rect 252388 298012 252394 298076
rect 252553 298074 252619 298077
rect 253606 298074 253612 298076
rect 252553 298072 253612 298074
rect 252553 298016 252558 298072
rect 252614 298016 253612 298072
rect 252553 298014 253612 298016
rect 252553 298011 252619 298014
rect 253606 298012 253612 298014
rect 253676 298012 253682 298076
rect 258030 298074 258090 298148
rect 258165 298074 258231 298077
rect 258030 298072 258231 298074
rect 258030 298016 258170 298072
rect 258226 298016 258231 298072
rect 258030 298014 258231 298016
rect 258165 298011 258231 298014
rect 259453 298076 259519 298077
rect 259453 298072 259500 298076
rect 259564 298074 259570 298076
rect 260189 298074 260255 298077
rect 260598 298074 260604 298076
rect 259453 298016 259458 298072
rect 259453 298012 259500 298016
rect 259564 298014 259610 298074
rect 260189 298072 260604 298074
rect 260189 298016 260194 298072
rect 260250 298016 260604 298072
rect 260189 298014 260604 298016
rect 259564 298012 259570 298014
rect 259453 298011 259519 298012
rect 260189 298011 260255 298014
rect 260598 298012 260604 298014
rect 260668 298012 260674 298076
rect 261109 298074 261175 298077
rect 261710 298074 261770 298148
rect 261109 298072 261770 298074
rect 261109 298016 261114 298072
rect 261170 298016 261770 298072
rect 261109 298014 261770 298016
rect 261109 298011 261175 298014
rect 263542 298012 263548 298076
rect 263612 298074 263618 298076
rect 263685 298074 263751 298077
rect 263612 298072 263751 298074
rect 263612 298016 263690 298072
rect 263746 298016 263751 298072
rect 263612 298014 263751 298016
rect 263612 298012 263618 298014
rect 263685 298011 263751 298014
rect 265065 298074 265131 298077
rect 265206 298074 265266 298148
rect 265065 298072 265266 298074
rect 265065 298016 265070 298072
rect 265126 298016 265266 298072
rect 265065 298014 265266 298016
rect 265341 298074 265407 298077
rect 266353 298076 266419 298077
rect 265934 298074 265940 298076
rect 265341 298072 265940 298074
rect 265341 298016 265346 298072
rect 265402 298016 265940 298072
rect 265341 298014 265940 298016
rect 265065 298011 265131 298014
rect 265341 298011 265407 298014
rect 265934 298012 265940 298014
rect 266004 298012 266010 298076
rect 266302 298074 266308 298076
rect 266262 298014 266308 298074
rect 266372 298072 266419 298076
rect 266414 298016 266419 298072
rect 266302 298012 266308 298014
rect 266372 298012 266419 298016
rect 266353 298011 266419 298012
rect 267825 298074 267891 298077
rect 269757 298076 269823 298077
rect 268694 298074 268700 298076
rect 267825 298072 268700 298074
rect 267825 298016 267830 298072
rect 267886 298016 268700 298072
rect 267825 298014 268700 298016
rect 267825 298011 267891 298014
rect 268694 298012 268700 298014
rect 268764 298012 268770 298076
rect 269757 298072 269804 298076
rect 269868 298074 269874 298076
rect 270493 298074 270559 298077
rect 270902 298074 270908 298076
rect 269757 298016 269762 298072
rect 269757 298012 269804 298016
rect 269868 298014 269914 298074
rect 270493 298072 270908 298074
rect 270493 298016 270498 298072
rect 270554 298016 270908 298072
rect 270493 298014 270908 298016
rect 269868 298012 269874 298014
rect 269757 298011 269823 298012
rect 270493 298011 270559 298014
rect 270902 298012 270908 298014
rect 270972 298012 270978 298076
rect 271873 298074 271939 298077
rect 272198 298074 272258 298148
rect 271873 298072 272258 298074
rect 271873 298016 271878 298072
rect 271934 298016 272258 298072
rect 271873 298014 272258 298016
rect 273253 298076 273319 298077
rect 273253 298072 273300 298076
rect 273364 298074 273370 298076
rect 274633 298074 274699 298077
rect 275694 298074 275754 298148
rect 276062 298077 276122 298148
rect 273253 298016 273258 298072
rect 271873 298011 271939 298014
rect 273253 298012 273300 298016
rect 273364 298014 273410 298074
rect 274633 298072 275754 298074
rect 274633 298016 274638 298072
rect 274694 298016 275754 298072
rect 274633 298014 275754 298016
rect 276013 298072 276122 298077
rect 276013 298016 276018 298072
rect 276074 298016 276122 298072
rect 276013 298014 276122 298016
rect 276749 298074 276815 298077
rect 276974 298074 276980 298076
rect 276749 298072 276980 298074
rect 276749 298016 276754 298072
rect 276810 298016 276980 298072
rect 276749 298014 276980 298016
rect 273364 298012 273370 298014
rect 273253 298011 273319 298012
rect 274633 298011 274699 298014
rect 276013 298011 276079 298014
rect 276749 298011 276815 298014
rect 276974 298012 276980 298014
rect 277044 298012 277050 298076
rect 277485 298074 277551 298077
rect 278446 298074 278452 298076
rect 277485 298072 278452 298074
rect 277485 298016 277490 298072
rect 277546 298016 278452 298072
rect 277485 298014 278452 298016
rect 277485 298011 277551 298014
rect 278446 298012 278452 298014
rect 278516 298012 278522 298076
rect 278773 298074 278839 298077
rect 278998 298074 279004 298076
rect 278773 298072 279004 298074
rect 278773 298016 278778 298072
rect 278834 298016 279004 298072
rect 278773 298014 279004 298016
rect 278773 298011 278839 298014
rect 278998 298012 279004 298014
rect 279068 298012 279074 298076
rect 280153 298074 280219 298077
rect 280838 298074 280844 298076
rect 280153 298072 280844 298074
rect 280153 298016 280158 298072
rect 280214 298016 280844 298072
rect 280153 298014 280844 298016
rect 280153 298011 280219 298014
rect 280838 298012 280844 298014
rect 280908 298012 280914 298076
rect 282913 298074 282979 298077
rect 283422 298074 283482 298148
rect 300902 298077 300962 298148
rect 315806 298077 315866 298148
rect 282913 298072 283482 298074
rect 282913 298016 282918 298072
rect 282974 298016 283482 298072
rect 282913 298014 283482 298016
rect 285949 298076 286015 298077
rect 285949 298072 285996 298076
rect 286060 298074 286066 298076
rect 287605 298074 287671 298077
rect 288198 298074 288204 298076
rect 285949 298016 285954 298072
rect 282913 298011 282979 298014
rect 285949 298012 285996 298016
rect 286060 298014 286106 298074
rect 287605 298072 288204 298074
rect 287605 298016 287610 298072
rect 287666 298016 288204 298072
rect 287605 298014 288204 298016
rect 286060 298012 286066 298014
rect 285949 298011 286015 298012
rect 287605 298011 287671 298014
rect 288198 298012 288204 298014
rect 288268 298012 288274 298076
rect 289997 298074 290063 298077
rect 290958 298074 290964 298076
rect 289997 298072 290964 298074
rect 289997 298016 290002 298072
rect 290058 298016 290964 298072
rect 289997 298014 290964 298016
rect 289997 298011 290063 298014
rect 290958 298012 290964 298014
rect 291028 298012 291034 298076
rect 292573 298074 292639 298077
rect 293350 298074 293356 298076
rect 292573 298072 293356 298074
rect 292573 298016 292578 298072
rect 292634 298016 293356 298072
rect 292573 298014 293356 298016
rect 292573 298011 292639 298014
rect 293350 298012 293356 298014
rect 293420 298012 293426 298076
rect 295333 298074 295399 298077
rect 298461 298076 298527 298077
rect 295926 298074 295932 298076
rect 295333 298072 295932 298074
rect 295333 298016 295338 298072
rect 295394 298016 295932 298072
rect 295333 298014 295932 298016
rect 295333 298011 295399 298014
rect 295926 298012 295932 298014
rect 295996 298012 296002 298076
rect 298461 298072 298508 298076
rect 298572 298074 298578 298076
rect 298461 298016 298466 298072
rect 298461 298012 298508 298016
rect 298572 298014 298618 298074
rect 300853 298072 300962 298077
rect 300853 298016 300858 298072
rect 300914 298016 300962 298072
rect 300853 298014 300962 298016
rect 302325 298074 302391 298077
rect 303470 298074 303476 298076
rect 302325 298072 303476 298074
rect 302325 298016 302330 298072
rect 302386 298016 303476 298072
rect 302325 298014 303476 298016
rect 298572 298012 298578 298014
rect 298461 298011 298527 298012
rect 300853 298011 300919 298014
rect 302325 298011 302391 298014
rect 303470 298012 303476 298014
rect 303540 298012 303546 298076
rect 305085 298074 305151 298077
rect 308581 298076 308647 298077
rect 310973 298076 311039 298077
rect 305862 298074 305868 298076
rect 305085 298072 305868 298074
rect 305085 298016 305090 298072
rect 305146 298016 305868 298072
rect 305085 298014 305868 298016
rect 305085 298011 305151 298014
rect 305862 298012 305868 298014
rect 305932 298012 305938 298076
rect 308581 298072 308628 298076
rect 308692 298074 308698 298076
rect 308581 298016 308586 298072
rect 308581 298012 308628 298016
rect 308692 298014 308738 298074
rect 310973 298072 311020 298076
rect 311084 298074 311090 298076
rect 313273 298074 313339 298077
rect 313406 298074 313412 298076
rect 310973 298016 310978 298072
rect 308692 298012 308698 298014
rect 310973 298012 311020 298016
rect 311084 298014 311130 298074
rect 313273 298072 313412 298074
rect 313273 298016 313278 298072
rect 313334 298016 313412 298072
rect 313273 298014 313412 298016
rect 311084 298012 311090 298014
rect 308581 298011 308647 298012
rect 310973 298011 311039 298012
rect 313273 298011 313339 298014
rect 313406 298012 313412 298014
rect 313476 298012 313482 298076
rect 315757 298072 315866 298077
rect 315757 298016 315762 298072
rect 315818 298016 315866 298072
rect 315757 298014 315866 298016
rect 317413 298074 317479 298077
rect 320909 298076 320975 298077
rect 318374 298074 318380 298076
rect 317413 298072 318380 298074
rect 317413 298016 317418 298072
rect 317474 298016 318380 298072
rect 317413 298014 318380 298016
rect 315757 298011 315823 298014
rect 317413 298011 317479 298014
rect 318374 298012 318380 298014
rect 318444 298012 318450 298076
rect 320909 298072 320956 298076
rect 321020 298074 321026 298076
rect 322933 298074 322999 298077
rect 323342 298074 323348 298076
rect 320909 298016 320914 298072
rect 320909 298012 320956 298016
rect 321020 298014 321066 298074
rect 322933 298072 323348 298074
rect 322933 298016 322938 298072
rect 322994 298016 323348 298072
rect 322933 298014 323348 298016
rect 321020 298012 321026 298014
rect 320909 298011 320975 298012
rect 322933 298011 322999 298014
rect 323342 298012 323348 298014
rect 323412 298012 323418 298076
rect 325693 298074 325759 298077
rect 325926 298074 325986 298148
rect 343173 298076 343239 298077
rect 343357 298076 343423 298077
rect 343173 298074 343220 298076
rect 325693 298072 325986 298074
rect 325693 298016 325698 298072
rect 325754 298016 325986 298072
rect 325693 298014 325986 298016
rect 343128 298072 343220 298074
rect 343128 298016 343178 298072
rect 343128 298014 343220 298016
rect 325693 298011 325759 298014
rect 343173 298012 343220 298014
rect 343284 298012 343290 298076
rect 343357 298072 343404 298076
rect 343468 298074 343474 298076
rect 343357 298016 343362 298072
rect 343357 298012 343404 298016
rect 343468 298014 343514 298074
rect 343468 298012 343474 298014
rect 343173 298011 343239 298012
rect 343357 298011 343423 298012
rect 96521 297938 96587 297941
rect 95742 297936 96587 297938
rect 95742 297880 96526 297936
rect 96582 297880 96587 297936
rect 95742 297878 96587 297880
rect 93412 297876 93418 297878
rect 93669 297875 93735 297878
rect 96521 297875 96587 297878
rect 98126 297876 98132 297940
rect 98196 297938 98202 297940
rect 99097 297938 99163 297941
rect 98196 297936 99163 297938
rect 98196 297880 99102 297936
rect 99158 297880 99163 297936
rect 98196 297878 99163 297880
rect 98196 297876 98202 297878
rect 99097 297875 99163 297878
rect 236494 297876 236500 297940
rect 236564 297938 236570 297940
rect 237281 297938 237347 297941
rect 248321 297940 248387 297941
rect 248270 297938 248276 297940
rect 236564 297936 237347 297938
rect 236564 297880 237286 297936
rect 237342 297880 237347 297936
rect 236564 297878 237347 297880
rect 248230 297878 248276 297938
rect 248340 297936 248387 297940
rect 248382 297880 248387 297936
rect 236564 297876 236570 297878
rect 237281 297875 237347 297878
rect 248270 297876 248276 297878
rect 248340 297876 248387 297880
rect 248321 297875 248387 297876
rect 263593 297938 263659 297941
rect 263910 297938 263916 297940
rect 263593 297936 263916 297938
rect 263593 297880 263598 297936
rect 263654 297880 263916 297936
rect 263593 297878 263916 297880
rect 263593 297875 263659 297878
rect 263910 297876 263916 297878
rect 263980 297876 263986 297940
rect 266445 297938 266511 297941
rect 267590 297938 267596 297940
rect 266445 297936 267596 297938
rect 266445 297880 266450 297936
rect 266506 297880 267596 297936
rect 266445 297878 267596 297880
rect 266445 297875 266511 297878
rect 267590 297876 267596 297878
rect 267660 297876 267666 297940
rect 268009 297938 268075 297941
rect 268326 297938 268332 297940
rect 268009 297936 268332 297938
rect 268009 297880 268014 297936
rect 268070 297880 268332 297936
rect 268009 297878 268332 297880
rect 268009 297875 268075 297878
rect 268326 297876 268332 297878
rect 268396 297876 268402 297940
rect 270585 297938 270651 297941
rect 271086 297938 271092 297940
rect 270585 297936 271092 297938
rect 270585 297880 270590 297936
rect 270646 297880 271092 297936
rect 270585 297878 271092 297880
rect 270585 297875 270651 297878
rect 271086 297876 271092 297878
rect 271156 297876 271162 297940
rect 273345 297938 273411 297941
rect 273478 297938 273484 297940
rect 273345 297936 273484 297938
rect 273345 297880 273350 297936
rect 273406 297880 273484 297936
rect 273345 297878 273484 297880
rect 273345 297875 273411 297878
rect 273478 297876 273484 297878
rect 273548 297876 273554 297940
rect 67766 297740 67772 297804
rect 67836 297802 67842 297804
rect 68829 297802 68895 297805
rect 67836 297800 68895 297802
rect 67836 297744 68834 297800
rect 68890 297744 68895 297800
rect 67836 297742 68895 297744
rect 67836 297740 67842 297742
rect 68829 297739 68895 297742
rect 76966 297740 76972 297804
rect 77036 297802 77042 297804
rect 77201 297802 77267 297805
rect 77036 297800 77267 297802
rect 77036 297744 77206 297800
rect 77262 297744 77267 297800
rect 77036 297742 77267 297744
rect 77036 297740 77042 297742
rect 77201 297739 77267 297742
rect 98494 297740 98500 297804
rect 98564 297802 98570 297804
rect 99281 297802 99347 297805
rect 98564 297800 99347 297802
rect 98564 297744 99286 297800
rect 99342 297744 99347 297800
rect 98564 297742 99347 297744
rect 98564 297740 98570 297742
rect 99281 297739 99347 297742
rect 219198 297740 219204 297804
rect 219268 297802 219274 297804
rect 240542 297802 240548 297804
rect 219268 297742 240548 297802
rect 219268 297740 219274 297742
rect 240542 297740 240548 297742
rect 240612 297740 240618 297804
rect 245510 297740 245516 297804
rect 245580 297802 245586 297804
rect 258349 297802 258415 297805
rect 245580 297800 258415 297802
rect 245580 297744 258354 297800
rect 258410 297744 258415 297800
rect 245580 297742 258415 297744
rect 245580 297740 245586 297742
rect 258349 297739 258415 297742
rect 273437 297802 273503 297805
rect 274398 297802 274404 297804
rect 273437 297800 274404 297802
rect 273437 297744 273442 297800
rect 273498 297744 274404 297800
rect 273437 297742 274404 297744
rect 273437 297739 273503 297742
rect 274398 297740 274404 297742
rect 274468 297740 274474 297804
rect 143390 297604 143396 297668
rect 143460 297666 143466 297668
rect 232446 297666 232452 297668
rect 143460 297606 232452 297666
rect 143460 297604 143466 297606
rect 232446 297604 232452 297606
rect 232516 297604 232522 297668
rect 242934 297604 242940 297668
rect 243004 297666 243010 297668
rect 258574 297666 258580 297668
rect 243004 297606 258580 297666
rect 243004 297604 243010 297606
rect 258574 297604 258580 297606
rect 258644 297604 258650 297668
rect 83590 297468 83596 297532
rect 83660 297530 83666 297532
rect 258942 297530 258948 297532
rect 83660 297470 258948 297530
rect 83660 297468 83666 297470
rect 258942 297468 258948 297470
rect 259012 297468 259018 297532
rect 70710 297332 70716 297396
rect 70780 297394 70786 297396
rect 70780 297334 238770 297394
rect 70780 297332 70786 297334
rect 238710 297258 238770 297334
rect 259494 297258 259500 297260
rect 238710 297198 259500 297258
rect 259494 297196 259500 297198
rect 259564 297196 259570 297260
rect 254526 297060 254532 297124
rect 254596 297122 254602 297124
rect 259126 297122 259132 297124
rect 254596 297062 259132 297122
rect 254596 297060 254602 297062
rect 259126 297060 259132 297062
rect 259196 297060 259202 297124
rect 256182 296924 256188 296988
rect 256252 296986 256258 296988
rect 256601 296986 256667 296989
rect 256252 296984 256667 296986
rect 256252 296928 256606 296984
rect 256662 296928 256667 296984
rect 256252 296926 256667 296928
rect 256252 296924 256258 296926
rect 256601 296923 256667 296926
rect 276657 296986 276723 296989
rect 278078 296986 278084 296988
rect 276657 296984 278084 296986
rect 276657 296928 276662 296984
rect 276718 296928 278084 296984
rect 276657 296926 278084 296928
rect 276657 296923 276723 296926
rect 278078 296924 278084 296926
rect 278148 296924 278154 296988
rect 103830 296788 103836 296852
rect 103900 296850 103906 296852
rect 104801 296850 104867 296853
rect 103900 296848 104867 296850
rect 103900 296792 104806 296848
rect 104862 296792 104867 296848
rect 103900 296790 104867 296792
rect 103900 296788 103906 296790
rect 104801 296787 104867 296790
rect 238702 296788 238708 296852
rect 238772 296850 238778 296852
rect 240041 296850 240107 296853
rect 238772 296848 240107 296850
rect 238772 296792 240046 296848
rect 240102 296792 240107 296848
rect 238772 296790 240107 296792
rect 238772 296788 238778 296790
rect 240041 296787 240107 296790
rect 255313 296850 255379 296853
rect 255814 296850 255820 296852
rect 255313 296848 255820 296850
rect 255313 296792 255318 296848
rect 255374 296792 255820 296848
rect 255313 296790 255820 296792
rect 255313 296787 255379 296790
rect 255814 296788 255820 296790
rect 255884 296788 255890 296852
rect 256693 296850 256759 296853
rect 256918 296850 256924 296852
rect 256693 296848 256924 296850
rect 256693 296792 256698 296848
rect 256754 296792 256924 296848
rect 256693 296790 256924 296792
rect 256693 296787 256759 296790
rect 256918 296788 256924 296790
rect 256988 296788 256994 296852
rect 258073 296850 258139 296853
rect 260925 296852 260991 296853
rect 258390 296850 258396 296852
rect 258073 296848 258396 296850
rect 258073 296792 258078 296848
rect 258134 296792 258396 296848
rect 258073 296790 258396 296792
rect 258073 296787 258139 296790
rect 258390 296788 258396 296790
rect 258460 296788 258466 296852
rect 260925 296848 260972 296852
rect 261036 296850 261042 296852
rect 262213 296850 262279 296853
rect 262806 296850 262812 296852
rect 260925 296792 260930 296848
rect 260925 296788 260972 296792
rect 261036 296790 261082 296850
rect 262213 296848 262812 296850
rect 262213 296792 262218 296848
rect 262274 296792 262812 296848
rect 262213 296790 262812 296792
rect 261036 296788 261042 296790
rect 260925 296787 260991 296788
rect 262213 296787 262279 296790
rect 262806 296788 262812 296790
rect 262876 296788 262882 296852
rect 258349 296036 258415 296037
rect 258349 296034 258396 296036
rect 258304 296032 258396 296034
rect 258304 295976 258354 296032
rect 258304 295974 258396 295976
rect 258349 295972 258396 295974
rect 258460 295972 258466 296036
rect 258349 295971 258415 295972
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 70301 239458 70367 239461
rect 259678 239458 259684 239460
rect 70301 239456 259684 239458
rect 70301 239400 70306 239456
rect 70362 239400 259684 239456
rect 70301 239398 259684 239400
rect 70301 239395 70367 239398
rect 259678 239396 259684 239398
rect 259748 239396 259754 239460
rect 583520 232236 584960 232476
rect 74349 230210 74415 230213
rect 262806 230210 262812 230212
rect 74349 230208 262812 230210
rect 74349 230152 74354 230208
rect 74410 230152 262812 230208
rect 74349 230150 262812 230152
rect 74349 230147 74415 230150
rect 262806 230148 262812 230150
rect 262876 230148 262882 230212
rect 66161 230074 66227 230077
rect 262438 230074 262444 230076
rect 66161 230072 262444 230074
rect 66161 230016 66166 230072
rect 66222 230016 262444 230072
rect 66161 230014 262444 230016
rect 66161 230011 66227 230014
rect 262438 230012 262444 230014
rect 262508 230012 262514 230076
rect 64781 229938 64847 229941
rect 262254 229938 262260 229940
rect 64781 229936 262260 229938
rect 64781 229880 64786 229936
rect 64842 229880 262260 229936
rect 64781 229878 262260 229880
rect 64781 229875 64847 229878
rect 262254 229876 262260 229878
rect 262324 229876 262330 229940
rect 38377 229802 38443 229805
rect 38377 229800 258090 229802
rect 38377 229744 38382 229800
rect 38438 229744 258090 229800
rect 38377 229742 258090 229744
rect 38377 229739 38443 229742
rect 258030 229666 258090 229742
rect 262622 229666 262628 229668
rect 258030 229606 262628 229666
rect 262622 229604 262628 229606
rect 262692 229604 262698 229668
rect 259361 229530 259427 229533
rect 259361 229528 259562 229530
rect 259361 229472 259366 229528
rect 259422 229472 259562 229528
rect 259361 229470 259562 229472
rect 259361 229467 259427 229470
rect 259502 229160 259562 229470
rect 110321 228986 110387 228989
rect 110278 228984 110387 228986
rect 110278 228928 110326 228984
rect 110382 228928 110387 228984
rect 110278 228923 110387 228928
rect 110278 228616 110338 228923
rect -960 227884 480 228124
rect 259913 228034 259979 228037
rect 259870 228032 259979 228034
rect 259870 227976 259918 228032
rect 259974 227976 259979 228032
rect 259870 227971 259979 227976
rect 259870 227528 259930 227971
rect 108481 226266 108547 226269
rect 259821 226266 259887 226269
rect 108481 226264 110154 226266
rect 108481 226208 108486 226264
rect 108542 226208 110154 226264
rect 108481 226206 110154 226208
rect 108481 226203 108547 226206
rect 110094 225896 110154 226206
rect 259821 226264 259930 226266
rect 259821 226208 259826 226264
rect 259882 226208 259930 226264
rect 259821 226203 259930 226208
rect 259870 225896 259930 226203
rect 263501 224634 263567 224637
rect 259870 224632 263567 224634
rect 259870 224576 263506 224632
rect 263562 224576 263567 224632
rect 259870 224574 263567 224576
rect 259870 224400 259930 224574
rect 263501 224571 263567 224574
rect 107653 223546 107719 223549
rect 107653 223544 110154 223546
rect 107653 223488 107658 223544
rect 107714 223488 110154 223544
rect 107653 223486 110154 223488
rect 107653 223483 107719 223486
rect 110094 223176 110154 223486
rect 262949 223138 263015 223141
rect 259870 223136 263015 223138
rect 259870 223080 262954 223136
rect 263010 223080 263015 223136
rect 259870 223078 263015 223080
rect 259870 222768 259930 223078
rect 262949 223075 263015 223078
rect 262857 221778 262923 221781
rect 259870 221776 262923 221778
rect 259870 221720 262862 221776
rect 262918 221720 262923 221776
rect 259870 221718 262923 221720
rect 259870 221136 259930 221718
rect 262857 221715 262923 221718
rect 109585 220486 109651 220489
rect 109585 220484 110124 220486
rect 109585 220428 109590 220484
rect 109646 220428 110124 220484
rect 109585 220426 110124 220428
rect 109585 220423 109651 220426
rect 262673 220282 262739 220285
rect 259870 220280 262739 220282
rect 259870 220224 262678 220280
rect 262734 220224 262739 220280
rect 259870 220222 262739 220224
rect 259870 219640 259930 220222
rect 262673 220219 262739 220222
rect 583520 218908 584960 219148
rect 259870 217970 259930 218008
rect 263501 217970 263567 217973
rect 259870 217968 263567 217970
rect 259870 217912 263506 217968
rect 263562 217912 263567 217968
rect 259870 217910 263567 217912
rect 263501 217907 263567 217910
rect 107653 217834 107719 217837
rect 107653 217832 110154 217834
rect 107653 217776 107658 217832
rect 107714 217776 110154 217832
rect 107653 217774 110154 217776
rect 107653 217771 107719 217774
rect 110094 217736 110154 217774
rect 263501 216474 263567 216477
rect 259870 216472 263567 216474
rect 259870 216416 263506 216472
rect 263562 216416 263567 216472
rect 259870 216414 263567 216416
rect 259870 216376 259930 216414
rect 263501 216411 263567 216414
rect 108573 215250 108639 215253
rect 262673 215250 262739 215253
rect 108573 215248 110154 215250
rect 108573 215192 108578 215248
rect 108634 215192 110154 215248
rect 108573 215190 110154 215192
rect 108573 215187 108639 215190
rect 110094 215152 110154 215190
rect 259870 215248 262739 215250
rect 259870 215192 262678 215248
rect 262734 215192 262739 215248
rect 259870 215190 262739 215192
rect -960 214828 480 215068
rect 259870 214744 259930 215190
rect 262673 215187 262739 215190
rect 263501 213618 263567 213621
rect 259870 213616 263567 213618
rect 259870 213560 263506 213616
rect 263562 213560 263567 213616
rect 259870 213558 263567 213560
rect 259870 213248 259930 213558
rect 263501 213555 263567 213558
rect 108665 212530 108731 212533
rect 108665 212528 110154 212530
rect 108665 212472 108670 212528
rect 108726 212472 110154 212528
rect 108665 212470 110154 212472
rect 108665 212467 108731 212470
rect 110094 212432 110154 212470
rect 261201 212258 261267 212261
rect 259870 212256 261267 212258
rect 259870 212200 261206 212256
rect 261262 212200 261267 212256
rect 259870 212198 261267 212200
rect 259870 211616 259930 212198
rect 261201 212195 261267 212198
rect 263501 210626 263567 210629
rect 259870 210624 263567 210626
rect 259870 210568 263506 210624
rect 263562 210568 263567 210624
rect 259870 210566 263567 210568
rect 259870 209984 259930 210566
rect 263501 210563 263567 210566
rect 109401 209674 109467 209677
rect 110094 209674 110154 209712
rect 109401 209672 110154 209674
rect 109401 209616 109406 209672
rect 109462 209616 110154 209672
rect 109401 209614 110154 209616
rect 109401 209611 109467 209614
rect 259729 209130 259795 209133
rect 259686 209128 259795 209130
rect 259686 209072 259734 209128
rect 259790 209072 259795 209128
rect 259686 209067 259795 209072
rect 259686 208488 259746 209067
rect 108757 206954 108823 206957
rect 110094 206954 110154 206992
rect 262581 206954 262647 206957
rect 108757 206952 110154 206954
rect 108757 206896 108762 206952
rect 108818 206896 110154 206952
rect 108757 206894 110154 206896
rect 259870 206952 262647 206954
rect 259870 206896 262586 206952
rect 262642 206896 262647 206952
rect 259870 206894 262647 206896
rect 108757 206891 108823 206894
rect 259870 206856 259930 206894
rect 262581 206891 262647 206894
rect 259637 205594 259703 205597
rect 259637 205592 259746 205594
rect 259637 205536 259642 205592
rect 259698 205536 259746 205592
rect 583520 205580 584960 205820
rect 259637 205531 259746 205536
rect 259686 205224 259746 205531
rect 109493 204914 109559 204917
rect 109493 204912 110154 204914
rect 109493 204856 109498 204912
rect 109554 204856 110154 204912
rect 109493 204854 110154 204856
rect 109493 204851 109559 204854
rect 110094 204272 110154 204854
rect 263501 203962 263567 203965
rect 259870 203960 263567 203962
rect 259870 203904 263506 203960
rect 263562 203904 263567 203960
rect 259870 203902 263567 203904
rect 259870 203728 259930 203902
rect 263501 203899 263567 203902
rect 259545 202738 259611 202741
rect 259502 202736 259611 202738
rect 259502 202680 259550 202736
rect 259606 202680 259611 202736
rect 259502 202675 259611 202680
rect 109309 202330 109375 202333
rect 109309 202328 110154 202330
rect 109309 202272 109314 202328
rect 109370 202272 110154 202328
rect 109309 202270 110154 202272
rect 109309 202267 109375 202270
rect -960 201772 480 202012
rect 110094 201688 110154 202270
rect 259502 202096 259562 202675
rect 262489 201106 262555 201109
rect 259870 201104 262555 201106
rect 259870 201048 262494 201104
rect 262550 201048 262555 201104
rect 259870 201046 262555 201048
rect 259870 200464 259930 201046
rect 262489 201043 262555 201046
rect 109217 199610 109283 199613
rect 109217 199608 110154 199610
rect 109217 199552 109222 199608
rect 109278 199552 110154 199608
rect 109217 199550 110154 199552
rect 109217 199547 109283 199550
rect 110094 198968 110154 199550
rect 260281 198862 260347 198865
rect 259900 198860 260347 198862
rect 259900 198804 260286 198860
rect 260342 198804 260347 198860
rect 259900 198802 260347 198804
rect 260281 198799 260347 198802
rect 259310 197508 259316 197572
rect 259380 197508 259386 197572
rect 259318 197336 259378 197508
rect 108849 196890 108915 196893
rect 108849 196888 110154 196890
rect 108849 196832 108854 196888
rect 108910 196832 110154 196888
rect 108849 196830 110154 196832
rect 108849 196827 108915 196830
rect 110094 196248 110154 196830
rect 262397 195938 262463 195941
rect 259870 195936 262463 195938
rect 259870 195880 262402 195936
rect 262458 195880 262463 195936
rect 259870 195878 262463 195880
rect 259870 195704 259930 195878
rect 262397 195875 262463 195878
rect 262806 194578 262812 194580
rect 259870 194518 262812 194578
rect 109125 194170 109191 194173
rect 109125 194168 110154 194170
rect 109125 194112 109130 194168
rect 109186 194112 110154 194168
rect 109125 194110 110154 194112
rect 109125 194107 109191 194110
rect 110094 193528 110154 194110
rect 259870 194072 259930 194518
rect 262806 194516 262812 194518
rect 262876 194516 262882 194580
rect 260189 192606 260255 192609
rect 259900 192604 260255 192606
rect 259900 192548 260194 192604
rect 260250 192548 260255 192604
rect 259900 192546 260255 192548
rect 260189 192543 260255 192546
rect 583520 192388 584960 192628
rect 259453 191586 259519 191589
rect 259453 191584 259562 191586
rect 259453 191528 259458 191584
rect 259514 191528 259562 191584
rect 259453 191523 259562 191528
rect 109033 191450 109099 191453
rect 109033 191448 110154 191450
rect 109033 191392 109038 191448
rect 109094 191392 110154 191448
rect 109033 191390 110154 191392
rect 109033 191387 109099 191390
rect 110094 190808 110154 191390
rect 259502 190944 259562 191523
rect 262213 189954 262279 189957
rect 259870 189952 262279 189954
rect 259870 189896 262218 189952
rect 262274 189896 262279 189952
rect 259870 189894 262279 189896
rect 259870 189312 259930 189894
rect 262213 189891 262279 189894
rect -960 188716 480 188956
rect 107653 188866 107719 188869
rect 107653 188864 110154 188866
rect 107653 188808 107658 188864
rect 107714 188808 110154 188864
rect 107653 188806 110154 188808
rect 107653 188803 107719 188806
rect 110094 188224 110154 188806
rect 260097 187710 260163 187713
rect 259900 187708 260163 187710
rect 259900 187652 260102 187708
rect 260158 187652 260163 187708
rect 259900 187650 260163 187652
rect 260097 187647 260163 187650
rect 259310 186356 259316 186420
rect 259380 186356 259386 186420
rect 259318 186184 259378 186356
rect 107653 186146 107719 186149
rect 107653 186144 110154 186146
rect 107653 186088 107658 186144
rect 107714 186088 110154 186144
rect 107653 186086 110154 186088
rect 107653 186083 107719 186086
rect 110094 185504 110154 186086
rect 259678 184860 259684 184924
rect 259748 184860 259754 184924
rect 259686 184552 259746 184860
rect 262622 183562 262628 183564
rect 259870 183502 262628 183562
rect 108941 183426 109007 183429
rect 108941 183424 110154 183426
rect 108941 183368 108946 183424
rect 109002 183368 110154 183424
rect 108941 183366 110154 183368
rect 108941 183363 109007 183366
rect 110094 182784 110154 183366
rect 259870 182920 259930 183502
rect 262622 183500 262628 183502
rect 262692 183500 262698 183564
rect 262305 182066 262371 182069
rect 259870 182064 262371 182066
rect 259870 182008 262310 182064
rect 262366 182008 262371 182064
rect 259870 182006 262371 182008
rect 259870 181424 259930 182006
rect 262305 182003 262371 182006
rect 107653 180706 107719 180709
rect 107653 180704 110154 180706
rect 107653 180648 107658 180704
rect 107714 180648 110154 180704
rect 107653 180646 110154 180648
rect 107653 180643 107719 180646
rect 110094 180064 110154 180646
rect 261109 180298 261175 180301
rect 259870 180296 261175 180298
rect 259870 180240 261114 180296
rect 261170 180240 261175 180296
rect 259870 180238 261175 180240
rect 259870 179792 259930 180238
rect 261109 180235 261175 180238
rect 583520 179060 584960 179300
rect 261017 178802 261083 178805
rect 259870 178800 261083 178802
rect 259870 178744 261022 178800
rect 261078 178744 261083 178800
rect 259870 178742 261083 178744
rect 259870 178160 259930 178742
rect 261017 178739 261083 178742
rect 107653 177986 107719 177989
rect 107653 177984 110154 177986
rect 107653 177928 107658 177984
rect 107714 177928 110154 177984
rect 107653 177926 110154 177928
rect 107653 177923 107719 177926
rect 110094 177344 110154 177926
rect 262438 177306 262444 177308
rect 259870 177246 262444 177306
rect 259870 176664 259930 177246
rect 262438 177244 262444 177246
rect 262508 177244 262514 177308
rect -960 175796 480 176036
rect 108389 175266 108455 175269
rect 108389 175264 110154 175266
rect 108389 175208 108394 175264
rect 108450 175208 110154 175264
rect 108389 175206 110154 175208
rect 108389 175203 108455 175206
rect 110094 174760 110154 175206
rect 259310 175204 259316 175268
rect 259380 175204 259386 175268
rect 259318 175032 259378 175204
rect 260925 173906 260991 173909
rect 259870 173904 260991 173906
rect 259870 173848 260930 173904
rect 260986 173848 260991 173904
rect 259870 173846 260991 173848
rect 259870 173400 259930 173846
rect 260925 173843 260991 173846
rect 107653 172410 107719 172413
rect 260005 172410 260071 172413
rect 107653 172408 110154 172410
rect 107653 172352 107658 172408
rect 107714 172352 110154 172408
rect 107653 172350 110154 172352
rect 107653 172347 107719 172350
rect 110094 172040 110154 172350
rect 259870 172408 260071 172410
rect 259870 172352 260010 172408
rect 260066 172352 260071 172408
rect 259870 172350 260071 172352
rect 259870 171768 259930 172350
rect 260005 172347 260071 172350
rect 259494 170716 259500 170780
rect 259564 170716 259570 170780
rect 259502 170272 259562 170716
rect 107653 169690 107719 169693
rect 107653 169688 110154 169690
rect 107653 169632 107658 169688
rect 107714 169632 110154 169688
rect 107653 169630 110154 169632
rect 107653 169627 107719 169630
rect 110094 169320 110154 169630
rect 260833 169282 260899 169285
rect 259870 169280 260899 169282
rect 259870 169224 260838 169280
rect 260894 169224 260899 169280
rect 259870 169222 260899 169224
rect 259870 168640 259930 169222
rect 260833 169219 260899 169222
rect 262254 167650 262260 167652
rect 259870 167590 262260 167650
rect 259870 167008 259930 167590
rect 262254 167588 262260 167590
rect 262324 167588 262330 167652
rect 108205 166970 108271 166973
rect 108205 166968 110154 166970
rect 108205 166912 108210 166968
rect 108266 166912 110154 166968
rect 108205 166910 110154 166912
rect 108205 166907 108271 166910
rect 110094 166600 110154 166910
rect 583520 165732 584960 165972
rect 259870 165341 259930 165512
rect 259870 165336 259979 165341
rect 259870 165280 259918 165336
rect 259974 165280 259979 165336
rect 259870 165278 259979 165280
rect 259913 165275 259979 165278
rect 259310 164188 259316 164252
rect 259380 164188 259386 164252
rect 107653 164114 107719 164117
rect 107653 164112 110154 164114
rect 107653 164056 107658 164112
rect 107714 164056 110154 164112
rect 107653 164054 110154 164056
rect 107653 164051 107719 164054
rect 110094 163880 110154 164054
rect 259318 163880 259378 164188
rect -960 162740 480 162980
rect 259821 162754 259887 162757
rect 259821 162752 259930 162754
rect 259821 162696 259826 162752
rect 259882 162696 259930 162752
rect 259821 162691 259930 162696
rect 259870 162248 259930 162691
rect 107653 161394 107719 161397
rect 107653 161392 110154 161394
rect 107653 161336 107658 161392
rect 107714 161336 110154 161392
rect 107653 161334 110154 161336
rect 107653 161331 107719 161334
rect 110094 161296 110154 161334
rect 263041 161122 263107 161125
rect 259870 161120 263107 161122
rect 259870 161064 263046 161120
rect 263102 161064 263107 161120
rect 259870 161062 263107 161064
rect 259870 160752 259930 161062
rect 263041 161059 263107 161062
rect 216765 160442 216831 160445
rect 217174 160442 217180 160444
rect 216765 160440 217180 160442
rect 216765 160384 216770 160440
rect 216826 160384 217180 160440
rect 216765 160382 217180 160384
rect 216765 160379 216831 160382
rect 217174 160380 217180 160382
rect 217244 160380 217250 160444
rect 218881 160442 218947 160445
rect 219198 160442 219204 160444
rect 218881 160440 219204 160442
rect 218881 160384 218886 160440
rect 218942 160384 219204 160440
rect 218881 160382 219204 160384
rect 218881 160379 218947 160382
rect 219198 160380 219204 160382
rect 219268 160380 219274 160444
rect 215845 158538 215911 158541
rect 244222 158538 244228 158540
rect 215845 158536 244228 158538
rect 215845 158480 215850 158536
rect 215906 158480 244228 158536
rect 215845 158478 244228 158480
rect 215845 158475 215911 158478
rect 244222 158476 244228 158478
rect 244292 158476 244298 158540
rect 220721 158402 220787 158405
rect 245694 158402 245700 158404
rect 220721 158400 245700 158402
rect 220721 158344 220726 158400
rect 220782 158344 245700 158400
rect 220721 158342 245700 158344
rect 220721 158339 220787 158342
rect 245694 158340 245700 158342
rect 245764 158340 245770 158404
rect 217542 158204 217548 158268
rect 217612 158266 217618 158268
rect 223665 158266 223731 158269
rect 217612 158264 223731 158266
rect 217612 158208 223670 158264
rect 223726 158208 223731 158264
rect 217612 158206 223731 158208
rect 217612 158204 217618 158206
rect 223665 158203 223731 158206
rect 232446 158204 232452 158268
rect 232516 158266 232522 158268
rect 258165 158266 258231 158269
rect 232516 158264 258231 158266
rect 232516 158208 258170 158264
rect 258226 158208 258231 158264
rect 232516 158206 258231 158208
rect 232516 158204 232522 158206
rect 258165 158203 258231 158206
rect 217358 158068 217364 158132
rect 217428 158130 217434 158132
rect 222285 158130 222351 158133
rect 217428 158128 222351 158130
rect 217428 158072 222290 158128
rect 222346 158072 222351 158128
rect 217428 158070 222351 158072
rect 217428 158068 217434 158070
rect 222285 158067 222351 158070
rect 228909 158130 228975 158133
rect 253422 158130 253428 158132
rect 228909 158128 253428 158130
rect 228909 158072 228914 158128
rect 228970 158072 253428 158128
rect 228909 158070 253428 158072
rect 228909 158067 228975 158070
rect 253422 158068 253428 158070
rect 253492 158068 253498 158132
rect 129958 157932 129964 157996
rect 130028 157994 130034 157996
rect 251909 157994 251975 157997
rect 130028 157992 251975 157994
rect 130028 157936 251914 157992
rect 251970 157936 251975 157992
rect 130028 157934 251975 157936
rect 130028 157932 130034 157934
rect 251909 157931 251975 157934
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 256693 119506 256759 119509
rect 342253 119506 342319 119509
rect 256693 119504 260084 119506
rect 256693 119448 256698 119504
rect 256754 119448 260084 119504
rect 256693 119446 260084 119448
rect 339940 119504 342319 119506
rect 339940 119448 342258 119504
rect 342314 119448 342319 119504
rect 339940 119446 342319 119448
rect 256693 119443 256759 119446
rect 342253 119443 342319 119446
rect 256693 118690 256759 118693
rect 342253 118690 342319 118693
rect 256693 118688 260084 118690
rect 256693 118632 256698 118688
rect 256754 118632 260084 118688
rect 256693 118630 260084 118632
rect 339940 118688 342319 118690
rect 339940 118632 342258 118688
rect 342314 118632 342319 118688
rect 339940 118630 342319 118632
rect 256693 118627 256759 118630
rect 342253 118627 342319 118630
rect 256785 117874 256851 117877
rect 342345 117874 342411 117877
rect 256785 117872 260084 117874
rect 256785 117816 256790 117872
rect 256846 117816 260084 117872
rect 256785 117814 260084 117816
rect 339940 117872 342411 117874
rect 339940 117816 342350 117872
rect 342406 117816 342411 117872
rect 339940 117814 342411 117816
rect 256785 117811 256851 117814
rect 342345 117811 342411 117814
rect 256693 117058 256759 117061
rect 342253 117058 342319 117061
rect 256693 117056 260084 117058
rect 256693 117000 256698 117056
rect 256754 117000 260084 117056
rect 256693 116998 260084 117000
rect 339940 117056 342319 117058
rect 339940 117000 342258 117056
rect 342314 117000 342319 117056
rect 339940 116998 342319 117000
rect 256693 116995 256759 116998
rect 342253 116995 342319 116998
rect 256785 116242 256851 116245
rect 342345 116242 342411 116245
rect 256785 116240 260084 116242
rect 256785 116184 256790 116240
rect 256846 116184 260084 116240
rect 256785 116182 260084 116184
rect 339940 116240 342411 116242
rect 339940 116184 342350 116240
rect 342406 116184 342411 116240
rect 339940 116182 342411 116184
rect 256785 116179 256851 116182
rect 342345 116179 342411 116182
rect 256693 115426 256759 115429
rect 342253 115426 342319 115429
rect 256693 115424 260084 115426
rect 256693 115368 256698 115424
rect 256754 115368 260084 115424
rect 256693 115366 260084 115368
rect 339940 115424 342319 115426
rect 339940 115368 342258 115424
rect 342314 115368 342319 115424
rect 339940 115366 342319 115368
rect 256693 115363 256759 115366
rect 342253 115363 342319 115366
rect 256785 114610 256851 114613
rect 342345 114610 342411 114613
rect 256785 114608 260084 114610
rect 256785 114552 256790 114608
rect 256846 114552 260084 114608
rect 256785 114550 260084 114552
rect 339940 114608 342411 114610
rect 339940 114552 342350 114608
rect 342406 114552 342411 114608
rect 339940 114550 342411 114552
rect 256785 114547 256851 114550
rect 342345 114547 342411 114550
rect 256693 113794 256759 113797
rect 342253 113794 342319 113797
rect 256693 113792 260084 113794
rect 256693 113736 256698 113792
rect 256754 113736 260084 113792
rect 256693 113734 260084 113736
rect 339940 113792 342319 113794
rect 339940 113736 342258 113792
rect 342314 113736 342319 113792
rect 339940 113734 342319 113736
rect 256693 113731 256759 113734
rect 342253 113731 342319 113734
rect 256693 113114 256759 113117
rect 342253 113114 342319 113117
rect 256693 113112 260084 113114
rect 256693 113056 256698 113112
rect 256754 113056 260084 113112
rect 256693 113054 260084 113056
rect 339940 113112 342319 113114
rect 339940 113056 342258 113112
rect 342314 113056 342319 113112
rect 339940 113054 342319 113056
rect 256693 113051 256759 113054
rect 342253 113051 342319 113054
rect 583520 112692 584960 112932
rect 256785 112298 256851 112301
rect 342345 112298 342411 112301
rect 256785 112296 260084 112298
rect 256785 112240 256790 112296
rect 256846 112240 260084 112296
rect 256785 112238 260084 112240
rect 339940 112296 342411 112298
rect 339940 112240 342350 112296
rect 342406 112240 342411 112296
rect 339940 112238 342411 112240
rect 256785 112235 256851 112238
rect 342345 112235 342411 112238
rect 256693 111482 256759 111485
rect 342253 111482 342319 111485
rect 256693 111480 260084 111482
rect 256693 111424 256698 111480
rect 256754 111424 260084 111480
rect 256693 111422 260084 111424
rect 339940 111480 342319 111482
rect 339940 111424 342258 111480
rect 342314 111424 342319 111480
rect 339940 111422 342319 111424
rect 256693 111419 256759 111422
rect 342253 111419 342319 111422
rect -960 110516 480 110756
rect 256785 110666 256851 110669
rect 342345 110666 342411 110669
rect 256785 110664 260084 110666
rect 256785 110608 256790 110664
rect 256846 110608 260084 110664
rect 256785 110606 260084 110608
rect 339940 110664 342411 110666
rect 339940 110608 342350 110664
rect 342406 110608 342411 110664
rect 339940 110606 342411 110608
rect 256785 110603 256851 110606
rect 342345 110603 342411 110606
rect 256693 109850 256759 109853
rect 342253 109850 342319 109853
rect 256693 109848 260084 109850
rect 256693 109792 256698 109848
rect 256754 109792 260084 109848
rect 256693 109790 260084 109792
rect 339940 109848 342319 109850
rect 339940 109792 342258 109848
rect 342314 109792 342319 109848
rect 339940 109790 342319 109792
rect 256693 109787 256759 109790
rect 342253 109787 342319 109790
rect 256693 109034 256759 109037
rect 342253 109034 342319 109037
rect 256693 109032 260084 109034
rect 256693 108976 256698 109032
rect 256754 108976 260084 109032
rect 256693 108974 260084 108976
rect 339940 109032 342319 109034
rect 339940 108976 342258 109032
rect 342314 108976 342319 109032
rect 339940 108974 342319 108976
rect 256693 108971 256759 108974
rect 342253 108971 342319 108974
rect 256785 108218 256851 108221
rect 342345 108218 342411 108221
rect 256785 108216 260084 108218
rect 256785 108160 256790 108216
rect 256846 108160 260084 108216
rect 256785 108158 260084 108160
rect 339940 108216 342411 108218
rect 339940 108160 342350 108216
rect 342406 108160 342411 108216
rect 339940 108158 342411 108160
rect 256785 108155 256851 108158
rect 342345 108155 342411 108158
rect 256693 107402 256759 107405
rect 342253 107402 342319 107405
rect 256693 107400 260084 107402
rect 256693 107344 256698 107400
rect 256754 107344 260084 107400
rect 256693 107342 260084 107344
rect 339940 107400 342319 107402
rect 339940 107344 342258 107400
rect 342314 107344 342319 107400
rect 339940 107342 342319 107344
rect 256693 107339 256759 107342
rect 342253 107339 342319 107342
rect 256785 106722 256851 106725
rect 342345 106722 342411 106725
rect 256785 106720 260084 106722
rect 256785 106664 256790 106720
rect 256846 106664 260084 106720
rect 256785 106662 260084 106664
rect 339940 106720 342411 106722
rect 339940 106664 342350 106720
rect 342406 106664 342411 106720
rect 339940 106662 342411 106664
rect 256785 106659 256851 106662
rect 342345 106659 342411 106662
rect 256693 105906 256759 105909
rect 342253 105906 342319 105909
rect 256693 105904 260084 105906
rect 256693 105848 256698 105904
rect 256754 105848 260084 105904
rect 256693 105846 260084 105848
rect 339940 105904 342319 105906
rect 339940 105848 342258 105904
rect 342314 105848 342319 105904
rect 339940 105846 342319 105848
rect 256693 105843 256759 105846
rect 342253 105843 342319 105846
rect 256785 105090 256851 105093
rect 342345 105090 342411 105093
rect 256785 105088 260084 105090
rect 256785 105032 256790 105088
rect 256846 105032 260084 105088
rect 256785 105030 260084 105032
rect 339940 105088 342411 105090
rect 339940 105032 342350 105088
rect 342406 105032 342411 105088
rect 339940 105030 342411 105032
rect 256785 105027 256851 105030
rect 342345 105027 342411 105030
rect 256693 104274 256759 104277
rect 342253 104274 342319 104277
rect 256693 104272 260084 104274
rect 256693 104216 256698 104272
rect 256754 104216 260084 104272
rect 256693 104214 260084 104216
rect 339940 104272 342319 104274
rect 339940 104216 342258 104272
rect 342314 104216 342319 104272
rect 339940 104214 342319 104216
rect 256693 104211 256759 104214
rect 342253 104211 342319 104214
rect 256693 103458 256759 103461
rect 342253 103458 342319 103461
rect 256693 103456 260084 103458
rect 256693 103400 256698 103456
rect 256754 103400 260084 103456
rect 256693 103398 260084 103400
rect 339940 103456 342319 103458
rect 339940 103400 342258 103456
rect 342314 103400 342319 103456
rect 339940 103398 342319 103400
rect 256693 103395 256759 103398
rect 342253 103395 342319 103398
rect 256785 102642 256851 102645
rect 342345 102642 342411 102645
rect 256785 102640 260084 102642
rect 256785 102584 256790 102640
rect 256846 102584 260084 102640
rect 256785 102582 260084 102584
rect 339940 102640 342411 102642
rect 339940 102584 342350 102640
rect 342406 102584 342411 102640
rect 339940 102582 342411 102584
rect 256785 102579 256851 102582
rect 342345 102579 342411 102582
rect 256693 101826 256759 101829
rect 342253 101826 342319 101829
rect 256693 101824 260084 101826
rect 256693 101768 256698 101824
rect 256754 101768 260084 101824
rect 256693 101766 260084 101768
rect 339940 101824 342319 101826
rect 339940 101768 342258 101824
rect 342314 101768 342319 101824
rect 339940 101766 342319 101768
rect 256693 101763 256759 101766
rect 342253 101763 342319 101766
rect 256785 101010 256851 101013
rect 342345 101010 342411 101013
rect 256785 101008 260084 101010
rect 256785 100952 256790 101008
rect 256846 100952 260084 101008
rect 256785 100950 260084 100952
rect 339940 101008 342411 101010
rect 339940 100952 342350 101008
rect 342406 100952 342411 101008
rect 339940 100950 342411 100952
rect 256785 100947 256851 100950
rect 342345 100947 342411 100950
rect 256693 100330 256759 100333
rect 342253 100330 342319 100333
rect 256693 100328 260084 100330
rect 256693 100272 256698 100328
rect 256754 100272 260084 100328
rect 256693 100270 260084 100272
rect 339940 100328 342319 100330
rect 339940 100272 342258 100328
rect 342314 100272 342319 100328
rect 339940 100270 342319 100272
rect 256693 100267 256759 100270
rect 342253 100267 342319 100270
rect 256785 99514 256851 99517
rect 342345 99514 342411 99517
rect 256785 99512 260084 99514
rect 256785 99456 256790 99512
rect 256846 99456 260084 99512
rect 256785 99454 260084 99456
rect 339940 99512 342411 99514
rect 339940 99456 342350 99512
rect 342406 99456 342411 99512
rect 339940 99454 342411 99456
rect 256785 99451 256851 99454
rect 342345 99451 342411 99454
rect 583520 99364 584960 99604
rect 256693 98698 256759 98701
rect 342253 98698 342319 98701
rect 256693 98696 260084 98698
rect 256693 98640 256698 98696
rect 256754 98640 260084 98696
rect 256693 98638 260084 98640
rect 339940 98696 342319 98698
rect 339940 98640 342258 98696
rect 342314 98640 342319 98696
rect 339940 98638 342319 98640
rect 256693 98635 256759 98638
rect 342253 98635 342319 98638
rect 256693 97882 256759 97885
rect 342253 97882 342319 97885
rect 256693 97880 260084 97882
rect 256693 97824 256698 97880
rect 256754 97824 260084 97880
rect 256693 97822 260084 97824
rect 339940 97880 342319 97882
rect 339940 97824 342258 97880
rect 342314 97824 342319 97880
rect 339940 97822 342319 97824
rect 256693 97819 256759 97822
rect 342253 97819 342319 97822
rect -960 97460 480 97700
rect 256785 97066 256851 97069
rect 342345 97066 342411 97069
rect 256785 97064 260084 97066
rect 256785 97008 256790 97064
rect 256846 97008 260084 97064
rect 256785 97006 260084 97008
rect 339940 97064 342411 97066
rect 339940 97008 342350 97064
rect 342406 97008 342411 97064
rect 339940 97006 342411 97008
rect 256785 97003 256851 97006
rect 342345 97003 342411 97006
rect 256693 96250 256759 96253
rect 342253 96250 342319 96253
rect 256693 96248 260084 96250
rect 256693 96192 256698 96248
rect 256754 96192 260084 96248
rect 256693 96190 260084 96192
rect 339940 96248 342319 96250
rect 339940 96192 342258 96248
rect 342314 96192 342319 96248
rect 339940 96190 342319 96192
rect 256693 96187 256759 96190
rect 342253 96187 342319 96190
rect 256785 95434 256851 95437
rect 342345 95434 342411 95437
rect 256785 95432 260084 95434
rect 256785 95376 256790 95432
rect 256846 95376 260084 95432
rect 256785 95374 260084 95376
rect 339940 95432 342411 95434
rect 339940 95376 342350 95432
rect 342406 95376 342411 95432
rect 339940 95374 342411 95376
rect 256785 95371 256851 95374
rect 342345 95371 342411 95374
rect 256693 94618 256759 94621
rect 342253 94618 342319 94621
rect 256693 94616 260084 94618
rect 256693 94560 256698 94616
rect 256754 94560 260084 94616
rect 256693 94558 260084 94560
rect 339940 94616 342319 94618
rect 339940 94560 342258 94616
rect 342314 94560 342319 94616
rect 339940 94558 342319 94560
rect 256693 94555 256759 94558
rect 342253 94555 342319 94558
rect 256693 93802 256759 93805
rect 342253 93802 342319 93805
rect 256693 93800 260084 93802
rect 256693 93744 256698 93800
rect 256754 93744 260084 93800
rect 256693 93742 260084 93744
rect 339940 93800 342319 93802
rect 339940 93744 342258 93800
rect 342314 93744 342319 93800
rect 339940 93742 342319 93744
rect 256693 93739 256759 93742
rect 342253 93739 342319 93742
rect 256785 93122 256851 93125
rect 342345 93122 342411 93125
rect 256785 93120 260084 93122
rect 256785 93064 256790 93120
rect 256846 93064 260084 93120
rect 256785 93062 260084 93064
rect 339940 93120 342411 93122
rect 339940 93064 342350 93120
rect 342406 93064 342411 93120
rect 339940 93062 342411 93064
rect 256785 93059 256851 93062
rect 342345 93059 342411 93062
rect 256693 92306 256759 92309
rect 342253 92306 342319 92309
rect 256693 92304 260084 92306
rect 256693 92248 256698 92304
rect 256754 92248 260084 92304
rect 256693 92246 260084 92248
rect 339940 92304 342319 92306
rect 339940 92248 342258 92304
rect 342314 92248 342319 92304
rect 339940 92246 342319 92248
rect 256693 92243 256759 92246
rect 342253 92243 342319 92246
rect 256785 91490 256851 91493
rect 342345 91490 342411 91493
rect 256785 91488 260084 91490
rect 256785 91432 256790 91488
rect 256846 91432 260084 91488
rect 256785 91430 260084 91432
rect 339940 91488 342411 91490
rect 339940 91432 342350 91488
rect 342406 91432 342411 91488
rect 339940 91430 342411 91432
rect 256785 91427 256851 91430
rect 342345 91427 342411 91430
rect 256693 90674 256759 90677
rect 342253 90674 342319 90677
rect 256693 90672 260084 90674
rect 256693 90616 256698 90672
rect 256754 90616 260084 90672
rect 256693 90614 260084 90616
rect 339940 90672 342319 90674
rect 339940 90616 342258 90672
rect 342314 90616 342319 90672
rect 339940 90614 342319 90616
rect 256693 90611 256759 90614
rect 342253 90611 342319 90614
rect 256785 89858 256851 89861
rect 342345 89858 342411 89861
rect 256785 89856 260084 89858
rect 256785 89800 256790 89856
rect 256846 89800 260084 89856
rect 256785 89798 260084 89800
rect 339940 89856 342411 89858
rect 339940 89800 342350 89856
rect 342406 89800 342411 89856
rect 339940 89798 342411 89800
rect 256785 89795 256851 89798
rect 342345 89795 342411 89798
rect 256693 89042 256759 89045
rect 342253 89042 342319 89045
rect 256693 89040 260084 89042
rect 256693 88984 256698 89040
rect 256754 88984 260084 89040
rect 256693 88982 260084 88984
rect 339940 89040 342319 89042
rect 339940 88984 342258 89040
rect 342314 88984 342319 89040
rect 339940 88982 342319 88984
rect 256693 88979 256759 88982
rect 342253 88979 342319 88982
rect 256693 88226 256759 88229
rect 342253 88226 342319 88229
rect 256693 88224 260084 88226
rect 256693 88168 256698 88224
rect 256754 88168 260084 88224
rect 256693 88166 260084 88168
rect 339940 88224 342319 88226
rect 339940 88168 342258 88224
rect 342314 88168 342319 88224
rect 339940 88166 342319 88168
rect 256693 88163 256759 88166
rect 342253 88163 342319 88166
rect 256785 87410 256851 87413
rect 342345 87410 342411 87413
rect 256785 87408 260084 87410
rect 256785 87352 256790 87408
rect 256846 87352 260084 87408
rect 256785 87350 260084 87352
rect 339940 87408 342411 87410
rect 339940 87352 342350 87408
rect 342406 87352 342411 87408
rect 339940 87350 342411 87352
rect 256785 87347 256851 87350
rect 342345 87347 342411 87350
rect 256693 86730 256759 86733
rect 342253 86730 342319 86733
rect 256693 86728 260084 86730
rect 256693 86672 256698 86728
rect 256754 86672 260084 86728
rect 256693 86670 260084 86672
rect 339940 86728 342319 86730
rect 339940 86672 342258 86728
rect 342314 86672 342319 86728
rect 339940 86670 342319 86672
rect 256693 86667 256759 86670
rect 342253 86667 342319 86670
rect 583520 86036 584960 86276
rect 256785 85914 256851 85917
rect 342345 85914 342411 85917
rect 256785 85912 260084 85914
rect 256785 85856 256790 85912
rect 256846 85856 260084 85912
rect 256785 85854 260084 85856
rect 339940 85912 342411 85914
rect 339940 85856 342350 85912
rect 342406 85856 342411 85912
rect 339940 85854 342411 85856
rect 256785 85851 256851 85854
rect 342345 85851 342411 85854
rect 256693 85098 256759 85101
rect 342253 85098 342319 85101
rect 256693 85096 260084 85098
rect 256693 85040 256698 85096
rect 256754 85040 260084 85096
rect 256693 85038 260084 85040
rect 339940 85096 342319 85098
rect 339940 85040 342258 85096
rect 342314 85040 342319 85096
rect 339940 85038 342319 85040
rect 256693 85035 256759 85038
rect 342253 85035 342319 85038
rect -960 84540 480 84780
rect 256785 84282 256851 84285
rect 342345 84282 342411 84285
rect 256785 84280 260084 84282
rect 256785 84224 256790 84280
rect 256846 84224 260084 84280
rect 256785 84222 260084 84224
rect 339940 84280 342411 84282
rect 339940 84224 342350 84280
rect 342406 84224 342411 84280
rect 339940 84222 342411 84224
rect 256785 84219 256851 84222
rect 342345 84219 342411 84222
rect 256693 83466 256759 83469
rect 342253 83466 342319 83469
rect 256693 83464 260084 83466
rect 256693 83408 256698 83464
rect 256754 83408 260084 83464
rect 256693 83406 260084 83408
rect 339940 83464 342319 83466
rect 339940 83408 342258 83464
rect 342314 83408 342319 83464
rect 339940 83406 342319 83408
rect 256693 83403 256759 83406
rect 342253 83403 342319 83406
rect 256693 82650 256759 82653
rect 342253 82650 342319 82653
rect 256693 82648 260084 82650
rect 256693 82592 256698 82648
rect 256754 82592 260084 82648
rect 256693 82590 260084 82592
rect 339940 82648 342319 82650
rect 339940 82592 342258 82648
rect 342314 82592 342319 82648
rect 339940 82590 342319 82592
rect 256693 82587 256759 82590
rect 342253 82587 342319 82590
rect 256785 81834 256851 81837
rect 342345 81834 342411 81837
rect 256785 81832 260084 81834
rect 256785 81776 256790 81832
rect 256846 81776 260084 81832
rect 256785 81774 260084 81776
rect 339940 81832 342411 81834
rect 339940 81776 342350 81832
rect 342406 81776 342411 81832
rect 339940 81774 342411 81776
rect 256785 81771 256851 81774
rect 342345 81771 342411 81774
rect 256693 81018 256759 81021
rect 342253 81018 342319 81021
rect 256693 81016 260084 81018
rect 256693 80960 256698 81016
rect 256754 80960 260084 81016
rect 256693 80958 260084 80960
rect 339940 81016 342319 81018
rect 339940 80960 342258 81016
rect 342314 80960 342319 81016
rect 339940 80958 342319 80960
rect 256693 80955 256759 80958
rect 342253 80955 342319 80958
rect 256785 80338 256851 80341
rect 342345 80338 342411 80341
rect 256785 80336 260084 80338
rect 256785 80280 256790 80336
rect 256846 80280 260084 80336
rect 256785 80278 260084 80280
rect 339940 80336 342411 80338
rect 339940 80280 342350 80336
rect 342406 80280 342411 80336
rect 339940 80278 342411 80280
rect 256785 80275 256851 80278
rect 342345 80275 342411 80278
rect 256693 79522 256759 79525
rect 342253 79522 342319 79525
rect 256693 79520 260084 79522
rect 256693 79464 256698 79520
rect 256754 79464 260084 79520
rect 256693 79462 260084 79464
rect 339940 79520 342319 79522
rect 339940 79464 342258 79520
rect 342314 79464 342319 79520
rect 339940 79462 342319 79464
rect 256693 79459 256759 79462
rect 342253 79459 342319 79462
rect 256785 78706 256851 78709
rect 342345 78706 342411 78709
rect 256785 78704 260084 78706
rect 256785 78648 256790 78704
rect 256846 78648 260084 78704
rect 256785 78646 260084 78648
rect 339940 78704 342411 78706
rect 339940 78648 342350 78704
rect 342406 78648 342411 78704
rect 339940 78646 342411 78648
rect 256785 78643 256851 78646
rect 342345 78643 342411 78646
rect 256693 77890 256759 77893
rect 342253 77890 342319 77893
rect 256693 77888 260084 77890
rect 256693 77832 256698 77888
rect 256754 77832 260084 77888
rect 256693 77830 260084 77832
rect 339940 77888 342319 77890
rect 339940 77832 342258 77888
rect 342314 77832 342319 77888
rect 339940 77830 342319 77832
rect 256693 77827 256759 77830
rect 342253 77827 342319 77830
rect 256693 77074 256759 77077
rect 342253 77074 342319 77077
rect 256693 77072 260084 77074
rect 256693 77016 256698 77072
rect 256754 77016 260084 77072
rect 256693 77014 260084 77016
rect 339940 77072 342319 77074
rect 339940 77016 342258 77072
rect 342314 77016 342319 77072
rect 339940 77014 342319 77016
rect 256693 77011 256759 77014
rect 342253 77011 342319 77014
rect 256785 76258 256851 76261
rect 342345 76258 342411 76261
rect 256785 76256 260084 76258
rect 256785 76200 256790 76256
rect 256846 76200 260084 76256
rect 256785 76198 260084 76200
rect 339940 76256 342411 76258
rect 339940 76200 342350 76256
rect 342406 76200 342411 76256
rect 339940 76198 342411 76200
rect 256785 76195 256851 76198
rect 342345 76195 342411 76198
rect 256693 75442 256759 75445
rect 342253 75442 342319 75445
rect 256693 75440 260084 75442
rect 256693 75384 256698 75440
rect 256754 75384 260084 75440
rect 256693 75382 260084 75384
rect 339940 75440 342319 75442
rect 339940 75384 342258 75440
rect 342314 75384 342319 75440
rect 339940 75382 342319 75384
rect 256693 75379 256759 75382
rect 342253 75379 342319 75382
rect 256785 74626 256851 74629
rect 342345 74626 342411 74629
rect 256785 74624 260084 74626
rect 256785 74568 256790 74624
rect 256846 74568 260084 74624
rect 256785 74566 260084 74568
rect 339940 74624 342411 74626
rect 339940 74568 342350 74624
rect 342406 74568 342411 74624
rect 339940 74566 342411 74568
rect 256785 74563 256851 74566
rect 342345 74563 342411 74566
rect 256693 73810 256759 73813
rect 342253 73810 342319 73813
rect 256693 73808 260084 73810
rect 256693 73752 256698 73808
rect 256754 73752 260084 73808
rect 256693 73750 260084 73752
rect 339940 73808 342319 73810
rect 339940 73752 342258 73808
rect 342314 73752 342319 73808
rect 339940 73750 342319 73752
rect 256693 73747 256759 73750
rect 342253 73747 342319 73750
rect 256693 73130 256759 73133
rect 342253 73130 342319 73133
rect 256693 73128 260084 73130
rect 256693 73072 256698 73128
rect 256754 73072 260084 73128
rect 256693 73070 260084 73072
rect 339940 73128 342319 73130
rect 339940 73072 342258 73128
rect 342314 73072 342319 73128
rect 339940 73070 342319 73072
rect 256693 73067 256759 73070
rect 342253 73067 342319 73070
rect 583520 72844 584960 73084
rect 256785 72314 256851 72317
rect 342345 72314 342411 72317
rect 256785 72312 260084 72314
rect 256785 72256 256790 72312
rect 256846 72256 260084 72312
rect 256785 72254 260084 72256
rect 339940 72312 342411 72314
rect 339940 72256 342350 72312
rect 342406 72256 342411 72312
rect 339940 72254 342411 72256
rect 256785 72251 256851 72254
rect 342345 72251 342411 72254
rect -960 71484 480 71724
rect 256693 71498 256759 71501
rect 342253 71498 342319 71501
rect 256693 71496 260084 71498
rect 256693 71440 256698 71496
rect 256754 71440 260084 71496
rect 256693 71438 260084 71440
rect 339940 71496 342319 71498
rect 339940 71440 342258 71496
rect 342314 71440 342319 71496
rect 339940 71438 342319 71440
rect 256693 71435 256759 71438
rect 342253 71435 342319 71438
rect 256785 70682 256851 70685
rect 342345 70682 342411 70685
rect 256785 70680 260084 70682
rect 256785 70624 256790 70680
rect 256846 70624 260084 70680
rect 256785 70622 260084 70624
rect 339940 70680 342411 70682
rect 339940 70624 342350 70680
rect 342406 70624 342411 70680
rect 339940 70622 342411 70624
rect 256785 70619 256851 70622
rect 342345 70619 342411 70622
rect 256693 69866 256759 69869
rect 342253 69866 342319 69869
rect 256693 69864 260084 69866
rect 256693 69808 256698 69864
rect 256754 69808 260084 69864
rect 256693 69806 260084 69808
rect 339940 69864 342319 69866
rect 339940 69808 342258 69864
rect 342314 69808 342319 69864
rect 339940 69806 342319 69808
rect 256693 69803 256759 69806
rect 342253 69803 342319 69806
rect 256785 69050 256851 69053
rect 342345 69050 342411 69053
rect 256785 69048 260084 69050
rect 256785 68992 256790 69048
rect 256846 68992 260084 69048
rect 256785 68990 260084 68992
rect 339940 69048 342411 69050
rect 339940 68992 342350 69048
rect 342406 68992 342411 69048
rect 339940 68990 342411 68992
rect 256785 68987 256851 68990
rect 342345 68987 342411 68990
rect 256693 68234 256759 68237
rect 342253 68234 342319 68237
rect 256693 68232 260084 68234
rect 256693 68176 256698 68232
rect 256754 68176 260084 68232
rect 256693 68174 260084 68176
rect 339940 68232 342319 68234
rect 339940 68176 342258 68232
rect 342314 68176 342319 68232
rect 339940 68174 342319 68176
rect 256693 68171 256759 68174
rect 342253 68171 342319 68174
rect 256693 67418 256759 67421
rect 342253 67418 342319 67421
rect 256693 67416 260084 67418
rect 256693 67360 256698 67416
rect 256754 67360 260084 67416
rect 256693 67358 260084 67360
rect 339940 67416 342319 67418
rect 339940 67360 342258 67416
rect 342314 67360 342319 67416
rect 339940 67358 342319 67360
rect 256693 67355 256759 67358
rect 342253 67355 342319 67358
rect 256785 66738 256851 66741
rect 342345 66738 342411 66741
rect 256785 66736 260084 66738
rect 256785 66680 256790 66736
rect 256846 66680 260084 66736
rect 256785 66678 260084 66680
rect 339940 66736 342411 66738
rect 339940 66680 342350 66736
rect 342406 66680 342411 66736
rect 339940 66678 342411 66680
rect 256785 66675 256851 66678
rect 342345 66675 342411 66678
rect 256693 65922 256759 65925
rect 342253 65922 342319 65925
rect 256693 65920 260084 65922
rect 256693 65864 256698 65920
rect 256754 65864 260084 65920
rect 256693 65862 260084 65864
rect 339940 65920 342319 65922
rect 339940 65864 342258 65920
rect 342314 65864 342319 65920
rect 339940 65862 342319 65864
rect 256693 65859 256759 65862
rect 342253 65859 342319 65862
rect 256785 65106 256851 65109
rect 342345 65106 342411 65109
rect 256785 65104 260084 65106
rect 256785 65048 256790 65104
rect 256846 65048 260084 65104
rect 256785 65046 260084 65048
rect 339940 65104 342411 65106
rect 339940 65048 342350 65104
rect 342406 65048 342411 65104
rect 339940 65046 342411 65048
rect 256785 65043 256851 65046
rect 342345 65043 342411 65046
rect 256693 64290 256759 64293
rect 342253 64290 342319 64293
rect 256693 64288 260084 64290
rect 256693 64232 256698 64288
rect 256754 64232 260084 64288
rect 256693 64230 260084 64232
rect 339940 64288 342319 64290
rect 339940 64232 342258 64288
rect 342314 64232 342319 64288
rect 339940 64230 342319 64232
rect 256693 64227 256759 64230
rect 342253 64227 342319 64230
rect 256693 63474 256759 63477
rect 342253 63474 342319 63477
rect 256693 63472 260084 63474
rect 256693 63416 256698 63472
rect 256754 63416 260084 63472
rect 256693 63414 260084 63416
rect 339940 63472 342319 63474
rect 339940 63416 342258 63472
rect 342314 63416 342319 63472
rect 339940 63414 342319 63416
rect 256693 63411 256759 63414
rect 342253 63411 342319 63414
rect 256785 62658 256851 62661
rect 342345 62658 342411 62661
rect 256785 62656 260084 62658
rect 256785 62600 256790 62656
rect 256846 62600 260084 62656
rect 256785 62598 260084 62600
rect 339940 62656 342411 62658
rect 339940 62600 342350 62656
rect 342406 62600 342411 62656
rect 339940 62598 342411 62600
rect 256785 62595 256851 62598
rect 342345 62595 342411 62598
rect 256693 61842 256759 61845
rect 342253 61842 342319 61845
rect 256693 61840 260084 61842
rect 256693 61784 256698 61840
rect 256754 61784 260084 61840
rect 256693 61782 260084 61784
rect 339940 61840 342319 61842
rect 339940 61784 342258 61840
rect 342314 61784 342319 61840
rect 339940 61782 342319 61784
rect 256693 61779 256759 61782
rect 342253 61779 342319 61782
rect 256785 61026 256851 61029
rect 342345 61026 342411 61029
rect 256785 61024 260084 61026
rect 256785 60968 256790 61024
rect 256846 60968 260084 61024
rect 256785 60966 260084 60968
rect 339940 61024 342411 61026
rect 339940 60968 342350 61024
rect 342406 60968 342411 61024
rect 339940 60966 342411 60968
rect 256785 60963 256851 60966
rect 342345 60963 342411 60966
rect 256693 60346 256759 60349
rect 342253 60346 342319 60349
rect 256693 60344 260084 60346
rect 256693 60288 256698 60344
rect 256754 60288 260084 60344
rect 256693 60286 260084 60288
rect 339940 60344 342319 60346
rect 339940 60288 342258 60344
rect 342314 60288 342319 60344
rect 339940 60286 342319 60288
rect 256693 60283 256759 60286
rect 342253 60283 342319 60286
rect 256785 59530 256851 59533
rect 342345 59530 342411 59533
rect 256785 59528 260084 59530
rect 256785 59472 256790 59528
rect 256846 59472 260084 59528
rect 256785 59470 260084 59472
rect 339940 59528 342411 59530
rect 339940 59472 342350 59528
rect 342406 59472 342411 59528
rect 583520 59516 584960 59756
rect 339940 59470 342411 59472
rect 256785 59467 256851 59470
rect 342345 59467 342411 59470
rect 256693 58714 256759 58717
rect 342253 58714 342319 58717
rect 256693 58712 260084 58714
rect -960 58428 480 58668
rect 256693 58656 256698 58712
rect 256754 58656 260084 58712
rect 256693 58654 260084 58656
rect 339940 58712 342319 58714
rect 339940 58656 342258 58712
rect 342314 58656 342319 58712
rect 339940 58654 342319 58656
rect 256693 58651 256759 58654
rect 342253 58651 342319 58654
rect 256693 57898 256759 57901
rect 342253 57898 342319 57901
rect 256693 57896 260084 57898
rect 256693 57840 256698 57896
rect 256754 57840 260084 57896
rect 256693 57838 260084 57840
rect 339940 57896 342319 57898
rect 339940 57840 342258 57896
rect 342314 57840 342319 57896
rect 339940 57838 342319 57840
rect 256693 57835 256759 57838
rect 342253 57835 342319 57838
rect 256785 57082 256851 57085
rect 342345 57082 342411 57085
rect 256785 57080 260084 57082
rect 256785 57024 256790 57080
rect 256846 57024 260084 57080
rect 256785 57022 260084 57024
rect 339940 57080 342411 57082
rect 339940 57024 342350 57080
rect 342406 57024 342411 57080
rect 339940 57022 342411 57024
rect 256785 57019 256851 57022
rect 342345 57019 342411 57022
rect 256693 56266 256759 56269
rect 342253 56266 342319 56269
rect 256693 56264 260084 56266
rect 256693 56208 256698 56264
rect 256754 56208 260084 56264
rect 256693 56206 260084 56208
rect 339940 56264 342319 56266
rect 339940 56208 342258 56264
rect 342314 56208 342319 56264
rect 339940 56206 342319 56208
rect 256693 56203 256759 56206
rect 342253 56203 342319 56206
rect 256785 55450 256851 55453
rect 342345 55450 342411 55453
rect 256785 55448 260084 55450
rect 256785 55392 256790 55448
rect 256846 55392 260084 55448
rect 256785 55390 260084 55392
rect 339940 55448 342411 55450
rect 339940 55392 342350 55448
rect 342406 55392 342411 55448
rect 339940 55390 342411 55392
rect 256785 55387 256851 55390
rect 342345 55387 342411 55390
rect 256693 54634 256759 54637
rect 342253 54634 342319 54637
rect 256693 54632 260084 54634
rect 256693 54576 256698 54632
rect 256754 54576 260084 54632
rect 256693 54574 260084 54576
rect 339940 54632 342319 54634
rect 339940 54576 342258 54632
rect 342314 54576 342319 54632
rect 339940 54574 342319 54576
rect 256693 54571 256759 54574
rect 342253 54571 342319 54574
rect 256693 53818 256759 53821
rect 342253 53818 342319 53821
rect 256693 53816 260084 53818
rect 256693 53760 256698 53816
rect 256754 53760 260084 53816
rect 256693 53758 260084 53760
rect 339940 53816 342319 53818
rect 339940 53760 342258 53816
rect 342314 53760 342319 53816
rect 339940 53758 342319 53760
rect 256693 53755 256759 53758
rect 342253 53755 342319 53758
rect 256785 53138 256851 53141
rect 342345 53138 342411 53141
rect 256785 53136 260084 53138
rect 256785 53080 256790 53136
rect 256846 53080 260084 53136
rect 256785 53078 260084 53080
rect 339940 53136 342411 53138
rect 339940 53080 342350 53136
rect 342406 53080 342411 53136
rect 339940 53078 342411 53080
rect 256785 53075 256851 53078
rect 342345 53075 342411 53078
rect 256693 52322 256759 52325
rect 342253 52322 342319 52325
rect 256693 52320 260084 52322
rect 256693 52264 256698 52320
rect 256754 52264 260084 52320
rect 256693 52262 260084 52264
rect 339940 52320 342319 52322
rect 339940 52264 342258 52320
rect 342314 52264 342319 52320
rect 339940 52262 342319 52264
rect 256693 52259 256759 52262
rect 342253 52259 342319 52262
rect 256785 51506 256851 51509
rect 342345 51506 342411 51509
rect 256785 51504 260084 51506
rect 256785 51448 256790 51504
rect 256846 51448 260084 51504
rect 256785 51446 260084 51448
rect 339940 51504 342411 51506
rect 339940 51448 342350 51504
rect 342406 51448 342411 51504
rect 339940 51446 342411 51448
rect 256785 51443 256851 51446
rect 342345 51443 342411 51446
rect 256693 50690 256759 50693
rect 342253 50690 342319 50693
rect 256693 50688 260084 50690
rect 256693 50632 256698 50688
rect 256754 50632 260084 50688
rect 256693 50630 260084 50632
rect 339940 50688 342319 50690
rect 339940 50632 342258 50688
rect 342314 50632 342319 50688
rect 339940 50630 342319 50632
rect 256693 50627 256759 50630
rect 342253 50627 342319 50630
rect 256785 49874 256851 49877
rect 342345 49874 342411 49877
rect 256785 49872 260084 49874
rect 256785 49816 256790 49872
rect 256846 49816 260084 49872
rect 256785 49814 260084 49816
rect 339940 49872 342411 49874
rect 339940 49816 342350 49872
rect 342406 49816 342411 49872
rect 339940 49814 342411 49816
rect 256785 49811 256851 49814
rect 342345 49811 342411 49814
rect 256693 49058 256759 49061
rect 342253 49058 342319 49061
rect 256693 49056 260084 49058
rect 256693 49000 256698 49056
rect 256754 49000 260084 49056
rect 256693 48998 260084 49000
rect 339940 49056 342319 49058
rect 339940 49000 342258 49056
rect 342314 49000 342319 49056
rect 339940 48998 342319 49000
rect 256693 48995 256759 48998
rect 342253 48995 342319 48998
rect 256693 48242 256759 48245
rect 342253 48242 342319 48245
rect 256693 48240 260084 48242
rect 256693 48184 256698 48240
rect 256754 48184 260084 48240
rect 256693 48182 260084 48184
rect 339940 48240 342319 48242
rect 339940 48184 342258 48240
rect 342314 48184 342319 48240
rect 339940 48182 342319 48184
rect 256693 48179 256759 48182
rect 342253 48179 342319 48182
rect 256785 47426 256851 47429
rect 342345 47426 342411 47429
rect 256785 47424 260084 47426
rect 256785 47368 256790 47424
rect 256846 47368 260084 47424
rect 256785 47366 260084 47368
rect 339940 47424 342411 47426
rect 339940 47368 342350 47424
rect 342406 47368 342411 47424
rect 339940 47366 342411 47368
rect 256785 47363 256851 47366
rect 342345 47363 342411 47366
rect 256693 46746 256759 46749
rect 342253 46746 342319 46749
rect 256693 46744 260084 46746
rect 256693 46688 256698 46744
rect 256754 46688 260084 46744
rect 256693 46686 260084 46688
rect 339940 46744 342319 46746
rect 339940 46688 342258 46744
rect 342314 46688 342319 46744
rect 339940 46686 342319 46688
rect 256693 46683 256759 46686
rect 342253 46683 342319 46686
rect 583520 46188 584960 46428
rect 256785 45930 256851 45933
rect 342345 45930 342411 45933
rect 256785 45928 260084 45930
rect 256785 45872 256790 45928
rect 256846 45872 260084 45928
rect 256785 45870 260084 45872
rect 339940 45928 342411 45930
rect 339940 45872 342350 45928
rect 342406 45872 342411 45928
rect 339940 45870 342411 45872
rect 256785 45867 256851 45870
rect 342345 45867 342411 45870
rect -960 45372 480 45612
rect 256693 45114 256759 45117
rect 342253 45114 342319 45117
rect 256693 45112 260084 45114
rect 256693 45056 256698 45112
rect 256754 45056 260084 45112
rect 256693 45054 260084 45056
rect 339940 45112 342319 45114
rect 339940 45056 342258 45112
rect 342314 45056 342319 45112
rect 339940 45054 342319 45056
rect 256693 45051 256759 45054
rect 342253 45051 342319 45054
rect 256785 44298 256851 44301
rect 342345 44298 342411 44301
rect 256785 44296 260084 44298
rect 256785 44240 256790 44296
rect 256846 44240 260084 44296
rect 256785 44238 260084 44240
rect 339940 44296 342411 44298
rect 339940 44240 342350 44296
rect 342406 44240 342411 44296
rect 339940 44238 342411 44240
rect 256785 44235 256851 44238
rect 342345 44235 342411 44238
rect 256693 43482 256759 43485
rect 342253 43482 342319 43485
rect 256693 43480 260084 43482
rect 256693 43424 256698 43480
rect 256754 43424 260084 43480
rect 256693 43422 260084 43424
rect 339940 43480 342319 43482
rect 339940 43424 342258 43480
rect 342314 43424 342319 43480
rect 339940 43422 342319 43424
rect 256693 43419 256759 43422
rect 342253 43419 342319 43422
rect 256693 42666 256759 42669
rect 342253 42666 342319 42669
rect 256693 42664 260084 42666
rect 256693 42608 256698 42664
rect 256754 42608 260084 42664
rect 256693 42606 260084 42608
rect 339940 42664 342319 42666
rect 339940 42608 342258 42664
rect 342314 42608 342319 42664
rect 339940 42606 342319 42608
rect 256693 42603 256759 42606
rect 342253 42603 342319 42606
rect 256785 41850 256851 41853
rect 342345 41850 342411 41853
rect 256785 41848 260084 41850
rect 256785 41792 256790 41848
rect 256846 41792 260084 41848
rect 256785 41790 260084 41792
rect 339940 41848 342411 41850
rect 339940 41792 342350 41848
rect 342406 41792 342411 41848
rect 339940 41790 342411 41792
rect 256785 41787 256851 41790
rect 342345 41787 342411 41790
rect 256693 41034 256759 41037
rect 342253 41034 342319 41037
rect 256693 41032 260084 41034
rect 256693 40976 256698 41032
rect 256754 40976 260084 41032
rect 256693 40974 260084 40976
rect 339940 41032 342319 41034
rect 339940 40976 342258 41032
rect 342314 40976 342319 41032
rect 339940 40974 342319 40976
rect 256693 40971 256759 40974
rect 342253 40971 342319 40974
rect 256785 40354 256851 40357
rect 342345 40354 342411 40357
rect 256785 40352 260084 40354
rect 256785 40296 256790 40352
rect 256846 40296 260084 40352
rect 256785 40294 260084 40296
rect 339940 40352 342411 40354
rect 339940 40296 342350 40352
rect 342406 40296 342411 40352
rect 339940 40294 342411 40296
rect 256785 40291 256851 40294
rect 342345 40291 342411 40294
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< via3 >>
rect 68692 386336 68756 386340
rect 68692 386280 68742 386336
rect 68742 386280 68756 386336
rect 68692 386276 68756 386280
rect 71084 386276 71148 386340
rect 78444 386336 78508 386340
rect 78444 386280 78494 386336
rect 78494 386280 78508 386336
rect 78444 386276 78508 386280
rect 88564 386276 88628 386340
rect 93532 386276 93596 386340
rect 96292 386276 96356 386340
rect 98500 386276 98564 386340
rect 100892 386276 100956 386340
rect 106044 386276 106108 386340
rect 108620 386276 108684 386340
rect 111012 386276 111076 386340
rect 115980 386276 116044 386340
rect 118556 386336 118620 386340
rect 118556 386280 118606 386336
rect 118606 386280 118620 386336
rect 118556 386276 118620 386280
rect 123524 386276 123588 386340
rect 125916 386276 125980 386340
rect 133644 386336 133708 386340
rect 133644 386280 133694 386336
rect 133694 386280 133708 386336
rect 133644 386276 133708 386280
rect 138428 386336 138492 386340
rect 138428 386280 138478 386336
rect 138478 386280 138492 386336
rect 138428 386276 138492 386280
rect 141004 386276 141068 386340
rect 143396 386336 143460 386340
rect 143396 386280 143446 386336
rect 143446 386280 143460 386336
rect 143396 386276 143460 386280
rect 158484 386336 158548 386340
rect 158484 386280 158534 386336
rect 158534 386280 158548 386336
rect 158484 386276 158548 386280
rect 159772 386336 159836 386340
rect 159772 386280 159822 386336
rect 159822 386280 159836 386336
rect 159772 386276 159836 386280
rect 248644 386276 248708 386340
rect 253428 386276 253492 386340
rect 256188 386276 256252 386340
rect 258396 386276 258460 386340
rect 260972 386276 261036 386340
rect 263548 386336 263612 386340
rect 263548 386280 263598 386336
rect 263598 386280 263612 386336
rect 263548 386276 263612 386280
rect 266124 386276 266188 386340
rect 268516 386276 268580 386340
rect 271092 386276 271156 386340
rect 273484 386276 273548 386340
rect 278452 386276 278516 386340
rect 280844 386276 280908 386340
rect 288572 386276 288636 386340
rect 295932 386276 295996 386340
rect 305868 386276 305932 386340
rect 311020 386276 311084 386340
rect 313596 386276 313660 386340
rect 318380 386276 318444 386340
rect 320956 386276 321020 386340
rect 323348 386276 323412 386340
rect 338436 386276 338500 386340
rect 339724 386276 339788 386340
rect 285996 386140 286060 386204
rect 290964 386140 291028 386204
rect 251036 386004 251100 386068
rect 316172 386004 316236 386068
rect 298508 385868 298572 385932
rect 303476 385868 303540 385932
rect 103652 385188 103716 385252
rect 73476 385052 73540 385116
rect 76236 385052 76300 385116
rect 81020 385112 81084 385116
rect 81020 385056 81070 385112
rect 81070 385056 81084 385112
rect 81020 385052 81084 385056
rect 83596 385112 83660 385116
rect 83596 385056 83646 385112
rect 83646 385056 83660 385112
rect 83596 385052 83660 385056
rect 86172 385052 86236 385116
rect 91140 385052 91204 385116
rect 113588 385052 113652 385116
rect 121132 385052 121196 385116
rect 128492 385052 128556 385116
rect 131068 385112 131132 385116
rect 131068 385056 131082 385112
rect 131082 385056 131132 385112
rect 131068 385052 131132 385056
rect 136036 385112 136100 385116
rect 136036 385056 136086 385112
rect 136086 385056 136100 385112
rect 136036 385052 136100 385056
rect 146156 385112 146220 385116
rect 146156 385056 146206 385112
rect 146206 385056 146220 385112
rect 146156 385052 146220 385056
rect 276060 385112 276124 385116
rect 276060 385056 276074 385112
rect 276074 385056 276124 385112
rect 276060 385052 276124 385056
rect 283604 385052 283668 385116
rect 293540 385052 293604 385116
rect 301084 385052 301148 385116
rect 308444 385052 308508 385116
rect 326108 385052 326172 385116
rect 350948 385112 351012 385116
rect 350948 385056 350998 385112
rect 350998 385056 351012 385112
rect 350948 385052 351012 385056
rect 170812 384160 170876 384164
rect 170812 384104 170862 384160
rect 170862 384104 170876 384160
rect 170812 384100 170876 384104
rect 217548 332692 217612 332756
rect 217364 330924 217428 330988
rect 217180 328068 217244 328132
rect 163222 299568 163286 299572
rect 163222 299512 163226 299568
rect 163226 299512 163282 299568
rect 163282 299512 163286 299568
rect 163222 299508 163286 299512
rect 163358 299568 163422 299572
rect 163358 299512 163410 299568
rect 163410 299512 163422 299568
rect 163358 299508 163422 299512
rect 55996 298148 56060 298212
rect 59676 298148 59740 298212
rect 63172 298148 63236 298212
rect 73660 298148 73724 298212
rect 85252 298148 85316 298212
rect 92244 298148 92308 298212
rect 95740 298148 95804 298212
rect 113404 298148 113468 298212
rect 120948 298148 121012 298212
rect 145972 298148 146036 298212
rect 258028 298148 258092 298212
rect 261708 298148 261772 298212
rect 265204 298148 265268 298212
rect 272196 298148 272260 298212
rect 275692 298148 275756 298212
rect 276060 298148 276124 298212
rect 283420 298148 283484 298212
rect 300900 298148 300964 298212
rect 315804 298148 315868 298212
rect 325924 298148 325988 298212
rect 57100 298012 57164 298076
rect 58204 298012 58268 298076
rect 60596 298072 60660 298076
rect 60596 298016 60646 298072
rect 60646 298016 60660 298072
rect 60596 298012 60660 298016
rect 61884 298012 61948 298076
rect 64276 298012 64340 298076
rect 65380 298012 65444 298076
rect 66484 298012 66548 298076
rect 68324 298012 68388 298076
rect 70164 298012 70228 298076
rect 71268 298012 71332 298076
rect 72372 298012 72436 298076
rect 74580 298012 74644 298076
rect 76052 298012 76116 298076
rect 78444 298072 78508 298076
rect 78444 298016 78494 298072
rect 78494 298016 78508 298072
rect 78444 298012 78508 298016
rect 79548 298012 79612 298076
rect 80652 298072 80716 298076
rect 80652 298016 80702 298072
rect 80702 298016 80716 298072
rect 80652 298012 80716 298016
rect 81020 298012 81084 298076
rect 81940 298012 82004 298076
rect 82860 298012 82924 298076
rect 83964 298072 84028 298076
rect 83964 298016 84014 298072
rect 84014 298016 84028 298072
rect 83964 298012 84028 298016
rect 85988 298012 86052 298076
rect 86356 298012 86420 298076
rect 88196 298072 88260 298076
rect 88196 298016 88210 298072
rect 88210 298016 88260 298072
rect 88196 298012 88260 298016
rect 88748 298012 88812 298076
rect 90956 298072 91020 298076
rect 90956 298016 91006 298072
rect 91006 298016 91020 298072
rect 90956 298012 91020 298016
rect 93532 298012 93596 298076
rect 94452 298012 94516 298076
rect 68692 297876 68756 297940
rect 73476 297876 73540 297940
rect 75868 297876 75932 297940
rect 78260 297876 78324 297940
rect 87644 297876 87708 297940
rect 89852 297876 89916 297940
rect 91140 297876 91204 297940
rect 93348 297876 93412 297940
rect 96292 298012 96356 298076
rect 97028 298012 97092 298076
rect 99052 298012 99116 298076
rect 100892 298012 100956 298076
rect 106044 298012 106108 298076
rect 108252 298012 108316 298076
rect 111012 298012 111076 298076
rect 115980 298072 116044 298076
rect 115980 298016 115994 298072
rect 115994 298016 116044 298072
rect 115980 298012 116044 298016
rect 118372 298012 118436 298076
rect 123524 298012 123588 298076
rect 125916 298072 125980 298076
rect 125916 298016 125930 298072
rect 125930 298016 125980 298072
rect 125916 298012 125980 298016
rect 128676 298012 128740 298076
rect 133460 298012 133524 298076
rect 136036 298072 136100 298076
rect 136036 298016 136086 298072
rect 136086 298016 136100 298072
rect 136036 298012 136100 298016
rect 138428 298012 138492 298076
rect 141004 298072 141068 298076
rect 141004 298016 141054 298072
rect 141054 298016 141068 298072
rect 141004 298012 141068 298016
rect 237052 298012 237116 298076
rect 238156 298072 238220 298076
rect 238156 298016 238170 298072
rect 238170 298016 238220 298072
rect 238156 298012 238220 298016
rect 241836 298012 241900 298076
rect 247724 298012 247788 298076
rect 248644 298012 248708 298076
rect 250116 298012 250180 298076
rect 250852 298012 250916 298076
rect 251220 298012 251284 298076
rect 252324 298012 252388 298076
rect 253612 298012 253676 298076
rect 259500 298072 259564 298076
rect 259500 298016 259514 298072
rect 259514 298016 259564 298072
rect 259500 298012 259564 298016
rect 260604 298012 260668 298076
rect 263548 298012 263612 298076
rect 265940 298012 266004 298076
rect 266308 298072 266372 298076
rect 266308 298016 266358 298072
rect 266358 298016 266372 298072
rect 266308 298012 266372 298016
rect 268700 298012 268764 298076
rect 269804 298072 269868 298076
rect 269804 298016 269818 298072
rect 269818 298016 269868 298072
rect 269804 298012 269868 298016
rect 270908 298012 270972 298076
rect 273300 298072 273364 298076
rect 273300 298016 273314 298072
rect 273314 298016 273364 298072
rect 273300 298012 273364 298016
rect 276980 298012 277044 298076
rect 278452 298012 278516 298076
rect 279004 298012 279068 298076
rect 280844 298012 280908 298076
rect 285996 298072 286060 298076
rect 285996 298016 286010 298072
rect 286010 298016 286060 298072
rect 285996 298012 286060 298016
rect 288204 298012 288268 298076
rect 290964 298012 291028 298076
rect 293356 298012 293420 298076
rect 295932 298012 295996 298076
rect 298508 298072 298572 298076
rect 298508 298016 298522 298072
rect 298522 298016 298572 298072
rect 298508 298012 298572 298016
rect 303476 298012 303540 298076
rect 305868 298012 305932 298076
rect 308628 298072 308692 298076
rect 308628 298016 308642 298072
rect 308642 298016 308692 298072
rect 308628 298012 308692 298016
rect 311020 298072 311084 298076
rect 311020 298016 311034 298072
rect 311034 298016 311084 298072
rect 311020 298012 311084 298016
rect 313412 298012 313476 298076
rect 318380 298012 318444 298076
rect 320956 298072 321020 298076
rect 320956 298016 320970 298072
rect 320970 298016 321020 298072
rect 320956 298012 321020 298016
rect 323348 298012 323412 298076
rect 343220 298072 343284 298076
rect 343220 298016 343234 298072
rect 343234 298016 343284 298072
rect 343220 298012 343284 298016
rect 343404 298072 343468 298076
rect 343404 298016 343418 298072
rect 343418 298016 343468 298072
rect 343404 298012 343468 298016
rect 98132 297876 98196 297940
rect 236500 297876 236564 297940
rect 248276 297936 248340 297940
rect 248276 297880 248326 297936
rect 248326 297880 248340 297936
rect 248276 297876 248340 297880
rect 263916 297876 263980 297940
rect 267596 297876 267660 297940
rect 268332 297876 268396 297940
rect 271092 297876 271156 297940
rect 273484 297876 273548 297940
rect 67772 297740 67836 297804
rect 76972 297740 77036 297804
rect 98500 297740 98564 297804
rect 219204 297740 219268 297804
rect 240548 297740 240612 297804
rect 245516 297740 245580 297804
rect 274404 297740 274468 297804
rect 143396 297604 143460 297668
rect 232452 297604 232516 297668
rect 242940 297604 243004 297668
rect 258580 297604 258644 297668
rect 83596 297468 83660 297532
rect 258948 297468 259012 297532
rect 70716 297332 70780 297396
rect 259500 297196 259564 297260
rect 254532 297060 254596 297124
rect 259132 297060 259196 297124
rect 256188 296924 256252 296988
rect 278084 296924 278148 296988
rect 103836 296788 103900 296852
rect 238708 296788 238772 296852
rect 255820 296788 255884 296852
rect 256924 296788 256988 296852
rect 258396 296788 258460 296852
rect 260972 296848 261036 296852
rect 260972 296792 260986 296848
rect 260986 296792 261036 296848
rect 260972 296788 261036 296792
rect 262812 296788 262876 296852
rect 258396 296032 258460 296036
rect 258396 295976 258410 296032
rect 258410 295976 258460 296032
rect 258396 295972 258460 295976
rect 259684 239396 259748 239460
rect 262812 230148 262876 230212
rect 262444 230012 262508 230076
rect 262260 229876 262324 229940
rect 262628 229604 262692 229668
rect 259316 197508 259380 197572
rect 262812 194516 262876 194580
rect 259316 186356 259380 186420
rect 259684 184860 259748 184924
rect 262628 183500 262692 183564
rect 262444 177244 262508 177308
rect 259316 175204 259380 175268
rect 259500 170716 259564 170780
rect 262260 167588 262324 167652
rect 259316 164188 259380 164252
rect 217180 160380 217244 160444
rect 219204 160380 219268 160444
rect 244228 158476 244292 158540
rect 245700 158340 245764 158404
rect 217548 158204 217612 158268
rect 232452 158204 232516 158268
rect 217364 158068 217428 158132
rect 253428 158068 253492 158132
rect 129964 157932 130028 157996
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 385308 38414 398898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 385308 42134 402618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 385308 45854 406338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 385308 49574 410058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 385308 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385308 60134 420618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 385308 63854 388338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 385308 67574 392058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 68691 386340 68757 386341
rect 68691 386276 68692 386340
rect 68756 386276 68757 386340
rect 68691 386275 68757 386276
rect 71083 386340 71149 386341
rect 71083 386276 71084 386340
rect 71148 386276 71149 386340
rect 71083 386275 71149 386276
rect 68694 383670 68754 386275
rect 71086 383670 71146 386275
rect 73794 385308 74414 398898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 385308 78134 402618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 78443 386340 78509 386341
rect 78443 386276 78444 386340
rect 78508 386276 78509 386340
rect 78443 386275 78509 386276
rect 73475 385116 73541 385117
rect 73475 385052 73476 385116
rect 73540 385052 73541 385116
rect 73475 385051 73541 385052
rect 76235 385116 76301 385117
rect 76235 385052 76236 385116
rect 76300 385052 76301 385116
rect 76235 385051 76301 385052
rect 73478 383670 73538 385051
rect 76238 383670 76298 385051
rect 68694 383610 68764 383670
rect 68704 383202 68764 383610
rect 71016 383610 71146 383670
rect 73464 383610 73538 383670
rect 76184 383610 76298 383670
rect 78446 383670 78506 386275
rect 81234 385308 81854 406338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 385308 85574 410058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 88563 386340 88629 386341
rect 88563 386276 88564 386340
rect 88628 386276 88629 386340
rect 88563 386275 88629 386276
rect 81019 385116 81085 385117
rect 81019 385052 81020 385116
rect 81084 385052 81085 385116
rect 81019 385051 81085 385052
rect 83595 385116 83661 385117
rect 83595 385052 83596 385116
rect 83660 385052 83661 385116
rect 83595 385051 83661 385052
rect 86171 385116 86237 385117
rect 86171 385052 86172 385116
rect 86236 385052 86237 385116
rect 86171 385051 86237 385052
rect 81022 383670 81082 385051
rect 83598 383670 83658 385051
rect 86174 383670 86234 385051
rect 88566 383670 88626 386275
rect 91794 385308 92414 416898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 93531 386340 93597 386341
rect 93531 386276 93532 386340
rect 93596 386276 93597 386340
rect 93531 386275 93597 386276
rect 91139 385116 91205 385117
rect 91139 385052 91140 385116
rect 91204 385052 91205 385116
rect 91139 385051 91205 385052
rect 78446 383610 78556 383670
rect 81022 383610 81140 383670
rect 71016 383202 71076 383610
rect 73464 383202 73524 383610
rect 76184 383202 76244 383610
rect 78496 383202 78556 383610
rect 81080 383202 81140 383610
rect 83528 383610 83658 383670
rect 86112 383610 86234 383670
rect 88560 383610 88626 383670
rect 91142 383670 91202 385051
rect 93534 383670 93594 386275
rect 95514 385308 96134 420618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 96291 386340 96357 386341
rect 96291 386276 96292 386340
rect 96356 386276 96357 386340
rect 96291 386275 96357 386276
rect 98499 386340 98565 386341
rect 98499 386276 98500 386340
rect 98564 386276 98565 386340
rect 98499 386275 98565 386276
rect 96294 383670 96354 386275
rect 98502 383670 98562 386275
rect 99234 385308 99854 388338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 100891 386340 100957 386341
rect 100891 386276 100892 386340
rect 100956 386276 100957 386340
rect 100891 386275 100957 386276
rect 91142 383610 91204 383670
rect 93534 383610 93652 383670
rect 83528 383202 83588 383610
rect 86112 383202 86172 383610
rect 88560 383202 88620 383610
rect 91144 383202 91204 383610
rect 93592 383202 93652 383610
rect 96176 383610 96354 383670
rect 98488 383610 98562 383670
rect 100894 383670 100954 386275
rect 102954 385308 103574 392058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 106043 386340 106109 386341
rect 106043 386276 106044 386340
rect 106108 386276 106109 386340
rect 106043 386275 106109 386276
rect 108619 386340 108685 386341
rect 108619 386276 108620 386340
rect 108684 386276 108685 386340
rect 108619 386275 108685 386276
rect 103651 385252 103717 385253
rect 103651 385188 103652 385252
rect 103716 385188 103717 385252
rect 103651 385187 103717 385188
rect 103654 383670 103714 385187
rect 106046 383670 106106 386275
rect 108622 383670 108682 386275
rect 109794 385308 110414 398898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 111011 386340 111077 386341
rect 111011 386276 111012 386340
rect 111076 386276 111077 386340
rect 111011 386275 111077 386276
rect 111014 383670 111074 386275
rect 113514 385308 114134 402618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 115979 386340 116045 386341
rect 115979 386276 115980 386340
rect 116044 386276 116045 386340
rect 115979 386275 116045 386276
rect 113587 385116 113653 385117
rect 113587 385052 113588 385116
rect 113652 385052 113653 385116
rect 113587 385051 113653 385052
rect 113590 383670 113650 385051
rect 115982 383670 116042 386275
rect 117234 385308 117854 406338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 502000 128414 524898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 502000 132134 528618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 502000 135854 532338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 502000 139574 536058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 502000 146414 506898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 502000 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 502000 153854 514338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 502000 157574 518058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 502000 164414 524898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 502000 168134 528618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 502000 171854 532338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 502000 175574 536058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 502000 182414 506898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 502000 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 502000 189854 514338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 502000 193574 518058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 502000 200414 524898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 502000 204134 528618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 502000 207854 532338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 502000 211574 536058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 502000 218414 506898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 502000 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 502000 225854 514338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 502000 229574 518058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 502000 236414 524898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 502000 240134 528618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 502000 243854 532338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 502000 247574 536058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 149568 489454 149888 489486
rect 149568 489218 149610 489454
rect 149846 489218 149888 489454
rect 149568 489134 149888 489218
rect 149568 488898 149610 489134
rect 149846 488898 149888 489134
rect 149568 488866 149888 488898
rect 180288 489454 180608 489486
rect 180288 489218 180330 489454
rect 180566 489218 180608 489454
rect 180288 489134 180608 489218
rect 180288 488898 180330 489134
rect 180566 488898 180608 489134
rect 180288 488866 180608 488898
rect 211008 489454 211328 489486
rect 211008 489218 211050 489454
rect 211286 489218 211328 489454
rect 211008 489134 211328 489218
rect 211008 488898 211050 489134
rect 211286 488898 211328 489134
rect 211008 488866 211328 488898
rect 241728 489454 242048 489486
rect 241728 489218 241770 489454
rect 242006 489218 242048 489454
rect 241728 489134 242048 489218
rect 241728 488898 241770 489134
rect 242006 488898 242048 489134
rect 241728 488866 242048 488898
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 134208 471454 134528 471486
rect 134208 471218 134250 471454
rect 134486 471218 134528 471454
rect 134208 471134 134528 471218
rect 134208 470898 134250 471134
rect 134486 470898 134528 471134
rect 134208 470866 134528 470898
rect 164928 471454 165248 471486
rect 164928 471218 164970 471454
rect 165206 471218 165248 471454
rect 164928 471134 165248 471218
rect 164928 470898 164970 471134
rect 165206 470898 165248 471134
rect 164928 470866 165248 470898
rect 195648 471454 195968 471486
rect 195648 471218 195690 471454
rect 195926 471218 195968 471454
rect 195648 471134 195968 471218
rect 195648 470898 195690 471134
rect 195926 470898 195968 471134
rect 195648 470866 195968 470898
rect 226368 471454 226688 471486
rect 226368 471218 226410 471454
rect 226646 471218 226688 471454
rect 226368 471134 226688 471218
rect 226368 470898 226410 471134
rect 226646 470898 226688 471134
rect 226368 470866 226688 470898
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 118555 386340 118621 386341
rect 118555 386276 118556 386340
rect 118620 386276 118621 386340
rect 118555 386275 118621 386276
rect 100894 383610 100996 383670
rect 103654 383610 103716 383670
rect 106046 383610 106164 383670
rect 96176 383202 96236 383610
rect 98488 383202 98548 383610
rect 100936 383202 100996 383610
rect 103656 383202 103716 383610
rect 106104 383202 106164 383610
rect 108552 383610 108682 383670
rect 111000 383610 111074 383670
rect 113584 383610 113650 383670
rect 115896 383610 116042 383670
rect 118558 383670 118618 386275
rect 120954 385308 121574 410058
rect 127794 453454 128414 458000
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 123523 386340 123589 386341
rect 123523 386276 123524 386340
rect 123588 386276 123589 386340
rect 123523 386275 123589 386276
rect 125915 386340 125981 386341
rect 125915 386276 125916 386340
rect 125980 386276 125981 386340
rect 125915 386275 125981 386276
rect 121131 385116 121197 385117
rect 121131 385052 121132 385116
rect 121196 385052 121197 385116
rect 121131 385051 121197 385052
rect 121134 383670 121194 385051
rect 123526 383670 123586 386275
rect 118558 383610 118676 383670
rect 108552 383202 108612 383610
rect 111000 383202 111060 383610
rect 113584 383202 113644 383610
rect 115896 383202 115956 383610
rect 118616 383202 118676 383610
rect 121064 383610 121194 383670
rect 123512 383610 123586 383670
rect 125918 383670 125978 386275
rect 127794 385308 128414 416898
rect 131514 457174 132134 458000
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385308 132134 420618
rect 135234 424894 135854 458000
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 133643 386340 133709 386341
rect 133643 386276 133644 386340
rect 133708 386276 133709 386340
rect 133643 386275 133709 386276
rect 128491 385116 128557 385117
rect 128491 385052 128492 385116
rect 128556 385052 128557 385116
rect 128491 385051 128557 385052
rect 131067 385116 131133 385117
rect 131067 385052 131068 385116
rect 131132 385052 131133 385116
rect 131067 385051 131133 385052
rect 128494 383670 128554 385051
rect 131070 383670 131130 385051
rect 133646 383670 133706 386275
rect 135234 385308 135854 388338
rect 138954 428614 139574 458000
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138427 386340 138493 386341
rect 138427 386276 138428 386340
rect 138492 386276 138493 386340
rect 138427 386275 138493 386276
rect 136035 385116 136101 385117
rect 136035 385052 136036 385116
rect 136100 385052 136101 385116
rect 136035 385051 136101 385052
rect 136038 383670 136098 385051
rect 125918 383610 126020 383670
rect 121064 383202 121124 383610
rect 123512 383202 123572 383610
rect 125960 383202 126020 383610
rect 128408 383610 128554 383670
rect 130992 383610 131130 383670
rect 133576 383610 133706 383670
rect 136024 383610 136098 383670
rect 138430 383670 138490 386275
rect 138954 385308 139574 392058
rect 145794 435454 146414 458000
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 141003 386340 141069 386341
rect 141003 386276 141004 386340
rect 141068 386276 141069 386340
rect 141003 386275 141069 386276
rect 143395 386340 143461 386341
rect 143395 386276 143396 386340
rect 143460 386276 143461 386340
rect 143395 386275 143461 386276
rect 141006 383670 141066 386275
rect 143398 383670 143458 386275
rect 145794 385308 146414 398898
rect 149514 439174 150134 458000
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 385308 150134 402618
rect 153234 442894 153854 458000
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 385308 153854 406338
rect 156954 446614 157574 458000
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 385308 157574 410058
rect 163794 453454 164414 458000
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 158483 386340 158549 386341
rect 158483 386276 158484 386340
rect 158548 386276 158549 386340
rect 158483 386275 158549 386276
rect 159771 386340 159837 386341
rect 159771 386276 159772 386340
rect 159836 386276 159837 386340
rect 159771 386275 159837 386276
rect 146155 385116 146221 385117
rect 146155 385052 146156 385116
rect 146220 385052 146221 385116
rect 146155 385051 146221 385052
rect 146158 383670 146218 385051
rect 158486 383670 158546 386275
rect 159774 383670 159834 386275
rect 163794 385308 164414 416898
rect 167514 457174 168134 458000
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385308 168134 420618
rect 171234 424894 171854 458000
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 385308 171854 388338
rect 174954 428614 175574 458000
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 385308 175574 392058
rect 181794 435454 182414 458000
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 170811 384164 170877 384165
rect 170811 384100 170812 384164
rect 170876 384100 170877 384164
rect 170811 384099 170877 384100
rect 138430 383610 138532 383670
rect 141006 383610 141116 383670
rect 128408 383202 128468 383610
rect 130992 383202 131052 383610
rect 133576 383202 133636 383610
rect 136024 383202 136084 383610
rect 138472 383202 138532 383610
rect 141056 383202 141116 383610
rect 143368 383610 143458 383670
rect 146088 383610 146218 383670
rect 158464 383610 158546 383670
rect 159688 383610 159834 383670
rect 170814 383670 170874 384099
rect 170814 383610 170900 383670
rect 143368 383202 143428 383610
rect 146088 383202 146148 383610
rect 158464 383202 158524 383610
rect 159688 383202 159748 383610
rect 170840 383202 170900 383610
rect 40272 381454 40620 381486
rect 40272 381218 40328 381454
rect 40564 381218 40620 381454
rect 40272 381134 40620 381218
rect 40272 380898 40328 381134
rect 40564 380898 40620 381134
rect 40272 380866 40620 380898
rect 176000 381454 176348 381486
rect 176000 381218 176056 381454
rect 176292 381218 176348 381454
rect 176000 381134 176348 381218
rect 176000 380898 176056 381134
rect 176292 380898 176348 381134
rect 176000 380866 176348 380898
rect 40952 363454 41300 363486
rect 40952 363218 41008 363454
rect 41244 363218 41300 363454
rect 40952 363134 41300 363218
rect 40952 362898 41008 363134
rect 41244 362898 41300 363134
rect 40952 362866 41300 362898
rect 175320 363454 175668 363486
rect 175320 363218 175376 363454
rect 175612 363218 175668 363454
rect 175320 363134 175668 363218
rect 175320 362898 175376 363134
rect 175612 362898 175668 363134
rect 175320 362866 175668 362898
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 40272 345454 40620 345486
rect 40272 345218 40328 345454
rect 40564 345218 40620 345454
rect 40272 345134 40620 345218
rect 40272 344898 40328 345134
rect 40564 344898 40620 345134
rect 40272 344866 40620 344898
rect 176000 345454 176348 345486
rect 176000 345218 176056 345454
rect 176292 345218 176348 345454
rect 176000 345134 176348 345218
rect 176000 344898 176056 345134
rect 176292 344898 176348 345134
rect 176000 344866 176348 344898
rect 40952 327454 41300 327486
rect 40952 327218 41008 327454
rect 41244 327218 41300 327454
rect 40952 327134 41300 327218
rect 40952 326898 41008 327134
rect 41244 326898 41300 327134
rect 40952 326866 41300 326898
rect 175320 327454 175668 327486
rect 175320 327218 175376 327454
rect 175612 327218 175668 327454
rect 175320 327134 175668 327218
rect 175320 326898 175376 327134
rect 175612 326898 175668 327134
rect 175320 326866 175668 326898
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 40272 309454 40620 309486
rect 40272 309218 40328 309454
rect 40564 309218 40620 309454
rect 40272 309134 40620 309218
rect 40272 308898 40328 309134
rect 40564 308898 40620 309134
rect 40272 308866 40620 308898
rect 176000 309454 176348 309486
rect 176000 309218 176056 309454
rect 176292 309218 176348 309454
rect 176000 309134 176348 309218
rect 176000 308898 176056 309134
rect 176292 308898 176348 309134
rect 176000 308866 176348 308898
rect 56056 299570 56116 300106
rect 57144 299570 57204 300106
rect 58232 299570 58292 300106
rect 55998 299510 56116 299570
rect 57102 299510 57204 299570
rect 58206 299510 58292 299570
rect 59592 299570 59652 300106
rect 60544 299570 60604 300106
rect 61768 299570 61828 300106
rect 63128 299570 63188 300106
rect 64216 299570 64276 300106
rect 65440 299570 65500 300106
rect 66528 299570 66588 300106
rect 59592 299510 59738 299570
rect 60544 299510 60658 299570
rect 61768 299510 61946 299570
rect 63128 299510 63234 299570
rect 64216 299510 64338 299570
rect 55998 298213 56058 299510
rect 55995 298212 56061 298213
rect 55995 298148 55996 298212
rect 56060 298148 56061 298212
rect 55995 298147 56061 298148
rect 57102 298077 57162 299510
rect 58206 298077 58266 299510
rect 59678 298213 59738 299510
rect 59675 298212 59741 298213
rect 59675 298148 59676 298212
rect 59740 298148 59741 298212
rect 59675 298147 59741 298148
rect 60598 298077 60658 299510
rect 61886 298077 61946 299510
rect 63174 298213 63234 299510
rect 63171 298212 63237 298213
rect 63171 298148 63172 298212
rect 63236 298148 63237 298212
rect 63171 298147 63237 298148
rect 64278 298077 64338 299510
rect 65382 299510 65500 299570
rect 66486 299510 66588 299570
rect 67616 299570 67676 300106
rect 68296 299570 68356 300106
rect 68704 299570 68764 300106
rect 67616 299510 67834 299570
rect 68296 299510 68386 299570
rect 65382 298077 65442 299510
rect 66486 298077 66546 299510
rect 57099 298076 57165 298077
rect 57099 298012 57100 298076
rect 57164 298012 57165 298076
rect 57099 298011 57165 298012
rect 58203 298076 58269 298077
rect 58203 298012 58204 298076
rect 58268 298012 58269 298076
rect 58203 298011 58269 298012
rect 60595 298076 60661 298077
rect 60595 298012 60596 298076
rect 60660 298012 60661 298076
rect 60595 298011 60661 298012
rect 61883 298076 61949 298077
rect 61883 298012 61884 298076
rect 61948 298012 61949 298076
rect 61883 298011 61949 298012
rect 64275 298076 64341 298077
rect 64275 298012 64276 298076
rect 64340 298012 64341 298076
rect 64275 298011 64341 298012
rect 65379 298076 65445 298077
rect 65379 298012 65380 298076
rect 65444 298012 65445 298076
rect 65379 298011 65445 298012
rect 66483 298076 66549 298077
rect 66483 298012 66484 298076
rect 66548 298012 66549 298076
rect 66483 298011 66549 298012
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 291454 38414 298000
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 295174 42134 298000
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 262894 45854 298000
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 266614 49574 298000
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 273454 56414 298000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 277174 60134 298000
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 280894 63854 298000
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 284614 67574 298000
rect 67774 297805 67834 299510
rect 68326 298077 68386 299510
rect 68694 299510 68764 299570
rect 70064 299570 70124 300106
rect 70744 299570 70804 300106
rect 71288 299570 71348 300106
rect 72376 299570 72436 300106
rect 70064 299510 70226 299570
rect 68323 298076 68389 298077
rect 68323 298012 68324 298076
rect 68388 298012 68389 298076
rect 68323 298011 68389 298012
rect 68694 297941 68754 299510
rect 70166 298077 70226 299510
rect 70718 299510 70804 299570
rect 71270 299510 71348 299570
rect 72374 299510 72436 299570
rect 73464 299570 73524 300106
rect 73600 299570 73660 300106
rect 74552 299570 74612 300106
rect 75912 299570 75972 300106
rect 73464 299510 73538 299570
rect 73600 299510 73722 299570
rect 74552 299510 74642 299570
rect 70163 298076 70229 298077
rect 70163 298012 70164 298076
rect 70228 298012 70229 298076
rect 70163 298011 70229 298012
rect 68691 297940 68757 297941
rect 68691 297876 68692 297940
rect 68756 297876 68757 297940
rect 68691 297875 68757 297876
rect 67771 297804 67837 297805
rect 67771 297740 67772 297804
rect 67836 297740 67837 297804
rect 67771 297739 67837 297740
rect 70718 297397 70778 299510
rect 71270 298077 71330 299510
rect 72374 298077 72434 299510
rect 71267 298076 71333 298077
rect 71267 298012 71268 298076
rect 71332 298012 71333 298076
rect 71267 298011 71333 298012
rect 72371 298076 72437 298077
rect 72371 298012 72372 298076
rect 72436 298012 72437 298076
rect 72371 298011 72437 298012
rect 73478 297941 73538 299510
rect 73662 298213 73722 299510
rect 73659 298212 73725 298213
rect 73659 298148 73660 298212
rect 73724 298148 73725 298212
rect 73659 298147 73725 298148
rect 74582 298077 74642 299510
rect 75870 299510 75972 299570
rect 76048 299570 76108 300106
rect 77000 299570 77060 300106
rect 76048 299510 76114 299570
rect 74579 298076 74645 298077
rect 74579 298012 74580 298076
rect 74644 298012 74645 298076
rect 74579 298011 74645 298012
rect 73475 297940 73541 297941
rect 73475 297876 73476 297940
rect 73540 297876 73541 297940
rect 73475 297875 73541 297876
rect 70715 297396 70781 297397
rect 70715 297332 70716 297396
rect 70780 297332 70781 297396
rect 70715 297331 70781 297332
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 291454 74414 298000
rect 75870 297941 75930 299510
rect 76054 298077 76114 299510
rect 76974 299510 77060 299570
rect 78088 299570 78148 300106
rect 78496 299570 78556 300106
rect 78088 299510 78322 299570
rect 76051 298076 76117 298077
rect 76051 298012 76052 298076
rect 76116 298012 76117 298076
rect 76051 298011 76117 298012
rect 75867 297940 75933 297941
rect 75867 297876 75868 297940
rect 75932 297876 75933 297940
rect 75867 297875 75933 297876
rect 76974 297805 77034 299510
rect 76971 297804 77037 297805
rect 76971 297740 76972 297804
rect 77036 297740 77037 297804
rect 76971 297739 77037 297740
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 295174 78134 298000
rect 78262 297941 78322 299510
rect 78446 299510 78556 299570
rect 79448 299570 79508 300106
rect 80672 299570 80732 300106
rect 81080 299570 81140 300106
rect 79448 299510 79610 299570
rect 78446 298077 78506 299510
rect 79550 298077 79610 299510
rect 80654 299510 80732 299570
rect 81022 299510 81140 299570
rect 81760 299570 81820 300106
rect 82848 299570 82908 300106
rect 83528 299570 83588 300106
rect 83936 299570 83996 300106
rect 85296 299570 85356 300106
rect 81760 299510 82002 299570
rect 82848 299510 82922 299570
rect 83528 299510 83658 299570
rect 83936 299510 84026 299570
rect 80654 298077 80714 299510
rect 81022 298077 81082 299510
rect 81942 298077 82002 299510
rect 82862 298077 82922 299510
rect 78443 298076 78509 298077
rect 78443 298012 78444 298076
rect 78508 298012 78509 298076
rect 78443 298011 78509 298012
rect 79547 298076 79613 298077
rect 79547 298012 79548 298076
rect 79612 298012 79613 298076
rect 79547 298011 79613 298012
rect 80651 298076 80717 298077
rect 80651 298012 80652 298076
rect 80716 298012 80717 298076
rect 80651 298011 80717 298012
rect 81019 298076 81085 298077
rect 81019 298012 81020 298076
rect 81084 298012 81085 298076
rect 81019 298011 81085 298012
rect 81939 298076 82005 298077
rect 81939 298012 81940 298076
rect 82004 298012 82005 298076
rect 81939 298011 82005 298012
rect 82859 298076 82925 298077
rect 82859 298012 82860 298076
rect 82924 298012 82925 298076
rect 82859 298011 82925 298012
rect 78259 297940 78325 297941
rect 78259 297876 78260 297940
rect 78324 297876 78325 297940
rect 78259 297875 78325 297876
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 262894 81854 298000
rect 83598 297533 83658 299510
rect 83966 298077 84026 299510
rect 85254 299510 85356 299570
rect 85976 299570 86036 300106
rect 86384 299570 86444 300106
rect 85976 299510 86050 299570
rect 85254 298213 85314 299510
rect 85251 298212 85317 298213
rect 85251 298148 85252 298212
rect 85316 298148 85317 298212
rect 85251 298147 85317 298148
rect 85990 298077 86050 299510
rect 86358 299510 86444 299570
rect 87608 299570 87668 300106
rect 88288 299570 88348 300106
rect 87608 299510 87706 299570
rect 86358 298077 86418 299510
rect 83963 298076 84029 298077
rect 83963 298012 83964 298076
rect 84028 298012 84029 298076
rect 83963 298011 84029 298012
rect 85987 298076 86053 298077
rect 85987 298012 85988 298076
rect 86052 298012 86053 298076
rect 85987 298011 86053 298012
rect 86355 298076 86421 298077
rect 86355 298012 86356 298076
rect 86420 298012 86421 298076
rect 86355 298011 86421 298012
rect 83595 297532 83661 297533
rect 83595 297468 83596 297532
rect 83660 297468 83661 297532
rect 83595 297467 83661 297468
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 266614 85574 298000
rect 87646 297941 87706 299510
rect 88198 299510 88348 299570
rect 88696 299570 88756 300106
rect 89784 299570 89844 300106
rect 91008 299570 91068 300106
rect 91144 299570 91204 300106
rect 88696 299510 88810 299570
rect 89784 299510 89914 299570
rect 88198 298077 88258 299510
rect 88750 298077 88810 299510
rect 88195 298076 88261 298077
rect 88195 298012 88196 298076
rect 88260 298012 88261 298076
rect 88195 298011 88261 298012
rect 88747 298076 88813 298077
rect 88747 298012 88748 298076
rect 88812 298012 88813 298076
rect 88747 298011 88813 298012
rect 89854 297941 89914 299510
rect 90958 299510 91068 299570
rect 91142 299510 91204 299570
rect 92232 299570 92292 300106
rect 93320 299570 93380 300106
rect 93592 299570 93652 300106
rect 92232 299510 92306 299570
rect 93320 299510 93410 299570
rect 90958 298077 91018 299510
rect 90955 298076 91021 298077
rect 90955 298012 90956 298076
rect 91020 298012 91021 298076
rect 90955 298011 91021 298012
rect 91142 297941 91202 299510
rect 92246 298213 92306 299510
rect 92243 298212 92309 298213
rect 92243 298148 92244 298212
rect 92308 298148 92309 298212
rect 92243 298147 92309 298148
rect 87643 297940 87709 297941
rect 87643 297876 87644 297940
rect 87708 297876 87709 297940
rect 87643 297875 87709 297876
rect 89851 297940 89917 297941
rect 89851 297876 89852 297940
rect 89916 297876 89917 297940
rect 89851 297875 89917 297876
rect 91139 297940 91205 297941
rect 91139 297876 91140 297940
rect 91204 297876 91205 297940
rect 91139 297875 91205 297876
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 273454 92414 298000
rect 93350 297941 93410 299510
rect 93534 299510 93652 299570
rect 94408 299570 94468 300106
rect 95768 299570 95828 300106
rect 94408 299510 94514 299570
rect 93534 298077 93594 299510
rect 94454 298077 94514 299510
rect 95742 299510 95828 299570
rect 96040 299570 96100 300106
rect 96992 299570 97052 300106
rect 98080 299570 98140 300106
rect 98488 299570 98548 300106
rect 99168 299570 99228 300106
rect 100936 299570 100996 300106
rect 96040 299510 96354 299570
rect 96992 299510 97090 299570
rect 98080 299510 98194 299570
rect 98488 299510 98562 299570
rect 95742 298213 95802 299510
rect 95739 298212 95805 298213
rect 95739 298148 95740 298212
rect 95804 298148 95805 298212
rect 95739 298147 95805 298148
rect 96294 298077 96354 299510
rect 97030 298077 97090 299510
rect 93531 298076 93597 298077
rect 93531 298012 93532 298076
rect 93596 298012 93597 298076
rect 93531 298011 93597 298012
rect 94451 298076 94517 298077
rect 94451 298012 94452 298076
rect 94516 298012 94517 298076
rect 94451 298011 94517 298012
rect 96291 298076 96357 298077
rect 96291 298012 96292 298076
rect 96356 298012 96357 298076
rect 96291 298011 96357 298012
rect 97027 298076 97093 298077
rect 97027 298012 97028 298076
rect 97092 298012 97093 298076
rect 97027 298011 97093 298012
rect 93347 297940 93413 297941
rect 93347 297876 93348 297940
rect 93412 297876 93413 297940
rect 93347 297875 93413 297876
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 277174 96134 298000
rect 98134 297941 98194 299510
rect 98131 297940 98197 297941
rect 98131 297876 98132 297940
rect 98196 297876 98197 297940
rect 98131 297875 98197 297876
rect 98502 297805 98562 299510
rect 99054 299510 99228 299570
rect 100894 299510 100996 299570
rect 103520 299570 103580 300106
rect 105968 299570 106028 300106
rect 108280 299570 108340 300106
rect 103520 299510 103714 299570
rect 105968 299510 106106 299570
rect 99054 298077 99114 299510
rect 100894 298077 100954 299510
rect 99051 298076 99117 298077
rect 99051 298012 99052 298076
rect 99116 298012 99117 298076
rect 99051 298011 99117 298012
rect 100891 298076 100957 298077
rect 100891 298012 100892 298076
rect 100956 298012 100957 298076
rect 100891 298011 100957 298012
rect 98499 297804 98565 297805
rect 98499 297740 98500 297804
rect 98564 297740 98565 297804
rect 98499 297739 98565 297740
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 280894 99854 298000
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 284614 103574 298000
rect 103654 296850 103714 299510
rect 106046 298077 106106 299510
rect 108254 299510 108340 299570
rect 111000 299570 111060 300106
rect 113448 299570 113508 300106
rect 111000 299510 111074 299570
rect 108254 298077 108314 299510
rect 111014 298077 111074 299510
rect 113406 299510 113508 299570
rect 115896 299570 115956 300106
rect 118480 299570 118540 300106
rect 115896 299510 116042 299570
rect 113406 298213 113466 299510
rect 113403 298212 113469 298213
rect 113403 298148 113404 298212
rect 113468 298148 113469 298212
rect 113403 298147 113469 298148
rect 115982 298077 116042 299510
rect 118374 299510 118540 299570
rect 120928 299570 120988 300106
rect 123512 299570 123572 300106
rect 125960 299570 126020 300106
rect 120928 299510 121010 299570
rect 123512 299510 123586 299570
rect 118374 298077 118434 299510
rect 120950 298213 121010 299510
rect 120947 298212 121013 298213
rect 120947 298148 120948 298212
rect 121012 298148 121013 298212
rect 120947 298147 121013 298148
rect 123526 298077 123586 299510
rect 125918 299510 126020 299570
rect 128544 299570 128604 300106
rect 130992 299570 131052 300106
rect 128544 299510 128738 299570
rect 125918 298077 125978 299510
rect 128678 298077 128738 299510
rect 130886 299510 131052 299570
rect 133440 299570 133500 300106
rect 135888 299570 135948 300106
rect 138472 299570 138532 300106
rect 133440 299510 133522 299570
rect 135888 299510 136098 299570
rect 106043 298076 106109 298077
rect 106043 298012 106044 298076
rect 106108 298012 106109 298076
rect 106043 298011 106109 298012
rect 108251 298076 108317 298077
rect 108251 298012 108252 298076
rect 108316 298012 108317 298076
rect 108251 298011 108317 298012
rect 111011 298076 111077 298077
rect 111011 298012 111012 298076
rect 111076 298012 111077 298076
rect 111011 298011 111077 298012
rect 115979 298076 116045 298077
rect 115979 298012 115980 298076
rect 116044 298012 116045 298076
rect 115979 298011 116045 298012
rect 118371 298076 118437 298077
rect 118371 298012 118372 298076
rect 118436 298012 118437 298076
rect 118371 298011 118437 298012
rect 123523 298076 123589 298077
rect 123523 298012 123524 298076
rect 123588 298012 123589 298076
rect 123523 298011 123589 298012
rect 125915 298076 125981 298077
rect 125915 298012 125916 298076
rect 125980 298012 125981 298076
rect 125915 298011 125981 298012
rect 128675 298076 128741 298077
rect 128675 298012 128676 298076
rect 128740 298012 128741 298076
rect 128675 298011 128741 298012
rect 103835 296852 103901 296853
rect 103835 296850 103836 296852
rect 103654 296790 103836 296850
rect 103835 296788 103836 296790
rect 103900 296788 103901 296852
rect 103835 296787 103901 296788
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 109794 291454 110414 298000
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 232000 110414 254898
rect 113514 295174 114134 298000
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 232000 114134 258618
rect 117234 262894 117854 298000
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 232000 117854 262338
rect 120954 266614 121574 298000
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 232000 121574 266058
rect 127794 273454 128414 298000
rect 130886 296730 130946 299510
rect 133462 298077 133522 299510
rect 136038 298077 136098 299510
rect 138430 299510 138532 299570
rect 140920 299570 140980 300106
rect 143368 299570 143428 300106
rect 145952 299570 146012 300106
rect 163224 299573 163284 300106
rect 163360 299573 163420 300106
rect 163221 299572 163287 299573
rect 140920 299510 141066 299570
rect 143368 299510 143458 299570
rect 145952 299510 146034 299570
rect 138430 298077 138490 299510
rect 141006 298077 141066 299510
rect 133459 298076 133525 298077
rect 133459 298012 133460 298076
rect 133524 298012 133525 298076
rect 133459 298011 133525 298012
rect 136035 298076 136101 298077
rect 136035 298012 136036 298076
rect 136100 298012 136101 298076
rect 136035 298011 136101 298012
rect 138427 298076 138493 298077
rect 138427 298012 138428 298076
rect 138492 298012 138493 298076
rect 138427 298011 138493 298012
rect 141003 298076 141069 298077
rect 141003 298012 141004 298076
rect 141068 298012 141069 298076
rect 141003 298011 141069 298012
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 232000 128414 236898
rect 129966 296670 130946 296730
rect 114208 219454 114528 219486
rect 114208 219218 114250 219454
rect 114486 219218 114528 219454
rect 114208 219134 114528 219218
rect 114208 218898 114250 219134
rect 114486 218898 114528 219134
rect 114208 218866 114528 218898
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 129568 201454 129888 201486
rect 129568 201218 129610 201454
rect 129846 201218 129888 201454
rect 129568 201134 129888 201218
rect 129568 200898 129610 201134
rect 129846 200898 129888 201134
rect 129568 200866 129888 200898
rect 114208 183454 114528 183486
rect 114208 183218 114250 183454
rect 114486 183218 114528 183454
rect 114208 183134 114528 183218
rect 114208 182898 114250 183134
rect 114486 182898 114528 183134
rect 114208 182866 114528 182898
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 129568 165454 129888 165486
rect 129568 165218 129610 165454
rect 129846 165218 129888 165454
rect 129568 165134 129888 165218
rect 129568 164898 129610 165134
rect 129846 164898 129888 165134
rect 129568 164866 129888 164898
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 147454 110414 158000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 151174 114134 158000
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 154894 117854 158000
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 122614 121574 158000
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 129454 128414 158000
rect 129966 157997 130026 296670
rect 131514 277174 132134 298000
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 232000 132134 240618
rect 135234 280894 135854 298000
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 232000 135854 244338
rect 138954 284614 139574 298000
rect 143398 297669 143458 299510
rect 145974 298213 146034 299510
rect 163221 299508 163222 299572
rect 163286 299508 163287 299572
rect 163221 299507 163287 299508
rect 163357 299572 163423 299573
rect 163357 299508 163358 299572
rect 163422 299508 163423 299572
rect 163357 299507 163423 299508
rect 145971 298212 146037 298213
rect 145971 298148 145972 298212
rect 146036 298148 146037 298212
rect 145971 298147 146037 298148
rect 143395 297668 143461 297669
rect 143395 297604 143396 297668
rect 143460 297604 143461 297668
rect 143395 297603 143461 297604
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 232000 139574 248058
rect 145794 291454 146414 298000
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 232000 146414 254898
rect 149514 295174 150134 298000
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 232000 150134 258618
rect 153234 262894 153854 298000
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 232000 153854 262338
rect 156954 266614 157574 298000
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 232000 157574 266058
rect 163794 273454 164414 298000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 232000 164414 236898
rect 167514 277174 168134 298000
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 232000 168134 240618
rect 171234 280894 171854 298000
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 232000 171854 244338
rect 174954 284614 175574 298000
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 232000 175574 248058
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 232000 182414 254898
rect 185514 439174 186134 458000
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 232000 186134 258618
rect 189234 442894 189854 458000
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 232000 189854 262338
rect 192954 446614 193574 458000
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 232000 193574 266058
rect 199794 453454 200414 458000
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 232000 200414 236898
rect 203514 457174 204134 458000
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 232000 204134 240618
rect 207234 424894 207854 458000
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 232000 207854 244338
rect 210954 428614 211574 458000
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 217794 435454 218414 458000
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 385308 218414 398898
rect 221514 439174 222134 458000
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 385308 222134 402618
rect 225234 442894 225854 458000
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 385308 225854 406338
rect 228954 446614 229574 458000
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 385308 229574 410058
rect 235794 453454 236414 458000
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 385308 236414 416898
rect 239514 457174 240134 458000
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385308 240134 420618
rect 243234 424894 243854 458000
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 385308 243854 388338
rect 246954 428614 247574 458000
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 385308 247574 392058
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 248643 386340 248709 386341
rect 248643 386276 248644 386340
rect 248708 386276 248709 386340
rect 248643 386275 248709 386276
rect 253427 386340 253493 386341
rect 253427 386276 253428 386340
rect 253492 386276 253493 386340
rect 253427 386275 253493 386276
rect 248646 383670 248706 386275
rect 251035 386068 251101 386069
rect 251035 386004 251036 386068
rect 251100 386004 251101 386068
rect 251035 386003 251101 386004
rect 251038 383670 251098 386003
rect 248646 383610 248764 383670
rect 248704 383202 248764 383610
rect 251016 383610 251098 383670
rect 253430 383670 253490 386275
rect 253794 385308 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 256187 386340 256253 386341
rect 256187 386276 256188 386340
rect 256252 386276 256253 386340
rect 256187 386275 256253 386276
rect 256190 383670 256250 386275
rect 257514 385308 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 258395 386340 258461 386341
rect 258395 386276 258396 386340
rect 258460 386276 258461 386340
rect 258395 386275 258461 386276
rect 260971 386340 261037 386341
rect 260971 386276 260972 386340
rect 261036 386276 261037 386340
rect 260971 386275 261037 386276
rect 253430 383610 253524 383670
rect 251016 383202 251076 383610
rect 253464 383202 253524 383610
rect 256184 383610 256250 383670
rect 258398 383670 258458 386275
rect 260974 383670 261034 386275
rect 261234 385308 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 263547 386340 263613 386341
rect 263547 386276 263548 386340
rect 263612 386276 263613 386340
rect 263547 386275 263613 386276
rect 263550 383670 263610 386275
rect 264954 385308 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 266123 386340 266189 386341
rect 266123 386276 266124 386340
rect 266188 386276 266189 386340
rect 266123 386275 266189 386276
rect 268515 386340 268581 386341
rect 268515 386276 268516 386340
rect 268580 386276 268581 386340
rect 268515 386275 268581 386276
rect 271091 386340 271157 386341
rect 271091 386276 271092 386340
rect 271156 386276 271157 386340
rect 271091 386275 271157 386276
rect 266126 383670 266186 386275
rect 258398 383610 258556 383670
rect 260974 383610 261140 383670
rect 256184 383202 256244 383610
rect 258496 383202 258556 383610
rect 261080 383202 261140 383610
rect 263528 383610 263610 383670
rect 266112 383610 266186 383670
rect 268518 383670 268578 386275
rect 271094 383670 271154 386275
rect 271794 385308 272414 416898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 273483 386340 273549 386341
rect 273483 386276 273484 386340
rect 273548 386276 273549 386340
rect 273483 386275 273549 386276
rect 273486 383670 273546 386275
rect 275514 385308 276134 420618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 278451 386340 278517 386341
rect 278451 386276 278452 386340
rect 278516 386276 278517 386340
rect 278451 386275 278517 386276
rect 276059 385116 276125 385117
rect 276059 385052 276060 385116
rect 276124 385052 276125 385116
rect 276059 385051 276125 385052
rect 276062 383670 276122 385051
rect 278454 383670 278514 386275
rect 279234 385308 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 280843 386340 280909 386341
rect 280843 386276 280844 386340
rect 280908 386276 280909 386340
rect 280843 386275 280909 386276
rect 280846 383670 280906 386275
rect 282954 385308 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 288571 386340 288637 386341
rect 288571 386276 288572 386340
rect 288636 386276 288637 386340
rect 288571 386275 288637 386276
rect 285995 386204 286061 386205
rect 285995 386140 285996 386204
rect 286060 386140 286061 386204
rect 285995 386139 286061 386140
rect 283603 385116 283669 385117
rect 283603 385052 283604 385116
rect 283668 385052 283669 385116
rect 283603 385051 283669 385052
rect 283606 383670 283666 385051
rect 285998 383670 286058 386139
rect 288574 383670 288634 386275
rect 289794 385308 290414 398898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 290963 386204 291029 386205
rect 290963 386140 290964 386204
rect 291028 386140 291029 386204
rect 290963 386139 291029 386140
rect 268518 383610 268620 383670
rect 271094 383610 271204 383670
rect 273486 383610 273652 383670
rect 276062 383610 276236 383670
rect 278454 383610 278548 383670
rect 280846 383610 280996 383670
rect 283606 383610 283716 383670
rect 285998 383610 286164 383670
rect 263528 383202 263588 383610
rect 266112 383202 266172 383610
rect 268560 383202 268620 383610
rect 271144 383202 271204 383610
rect 273592 383202 273652 383610
rect 276176 383202 276236 383610
rect 278488 383202 278548 383610
rect 280936 383202 280996 383610
rect 283656 383202 283716 383610
rect 286104 383202 286164 383610
rect 288552 383610 288634 383670
rect 290966 383670 291026 386139
rect 293514 385308 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 295931 386340 295997 386341
rect 295931 386276 295932 386340
rect 295996 386276 295997 386340
rect 295931 386275 295997 386276
rect 293539 385116 293605 385117
rect 293539 385052 293540 385116
rect 293604 385052 293605 385116
rect 293539 385051 293605 385052
rect 293542 383670 293602 385051
rect 295934 383670 295994 386275
rect 297234 385308 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 298507 385932 298573 385933
rect 298507 385868 298508 385932
rect 298572 385868 298573 385932
rect 298507 385867 298573 385868
rect 290966 383610 291060 383670
rect 293542 383610 293644 383670
rect 288552 383202 288612 383610
rect 291000 383202 291060 383610
rect 293584 383202 293644 383610
rect 295896 383610 295994 383670
rect 298510 383670 298570 385867
rect 300954 385308 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 305867 386340 305933 386341
rect 305867 386276 305868 386340
rect 305932 386276 305933 386340
rect 305867 386275 305933 386276
rect 303475 385932 303541 385933
rect 303475 385868 303476 385932
rect 303540 385868 303541 385932
rect 303475 385867 303541 385868
rect 301083 385116 301149 385117
rect 301083 385052 301084 385116
rect 301148 385052 301149 385116
rect 301083 385051 301149 385052
rect 301086 383670 301146 385051
rect 298510 383610 298676 383670
rect 295896 383202 295956 383610
rect 298616 383202 298676 383610
rect 301064 383610 301146 383670
rect 303478 383670 303538 385867
rect 305870 383670 305930 386275
rect 307794 385308 308414 416898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311019 386340 311085 386341
rect 311019 386276 311020 386340
rect 311084 386276 311085 386340
rect 311019 386275 311085 386276
rect 308443 385116 308509 385117
rect 308443 385052 308444 385116
rect 308508 385052 308509 385116
rect 308443 385051 308509 385052
rect 308446 383670 308506 385051
rect 311022 383670 311082 386275
rect 311514 385308 312134 420618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 313595 386340 313661 386341
rect 313595 386276 313596 386340
rect 313660 386276 313661 386340
rect 313595 386275 313661 386276
rect 313598 383670 313658 386275
rect 315234 385308 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318379 386340 318445 386341
rect 318379 386276 318380 386340
rect 318444 386276 318445 386340
rect 318379 386275 318445 386276
rect 316171 386068 316237 386069
rect 316171 386004 316172 386068
rect 316236 386004 316237 386068
rect 316171 386003 316237 386004
rect 316174 383670 316234 386003
rect 303478 383610 303572 383670
rect 305870 383610 306020 383670
rect 301064 383202 301124 383610
rect 303512 383202 303572 383610
rect 305960 383202 306020 383610
rect 308408 383610 308506 383670
rect 310992 383610 311082 383670
rect 313576 383610 313658 383670
rect 316024 383610 316234 383670
rect 318382 383670 318442 386275
rect 318954 385308 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 320955 386340 321021 386341
rect 320955 386276 320956 386340
rect 321020 386276 321021 386340
rect 320955 386275 321021 386276
rect 323347 386340 323413 386341
rect 323347 386276 323348 386340
rect 323412 386276 323413 386340
rect 323347 386275 323413 386276
rect 320958 383670 321018 386275
rect 323350 383670 323410 386275
rect 325794 385308 326414 398898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 385308 330134 402618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 385308 333854 406338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 385308 337574 410058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 338435 386340 338501 386341
rect 338435 386276 338436 386340
rect 338500 386276 338501 386340
rect 338435 386275 338501 386276
rect 339723 386340 339789 386341
rect 339723 386276 339724 386340
rect 339788 386276 339789 386340
rect 339723 386275 339789 386276
rect 326107 385116 326173 385117
rect 326107 385052 326108 385116
rect 326172 385052 326173 385116
rect 326107 385051 326173 385052
rect 326110 383670 326170 385051
rect 318382 383610 318532 383670
rect 320958 383610 321116 383670
rect 323350 383610 323428 383670
rect 308408 383202 308468 383610
rect 310992 383202 311052 383610
rect 313576 383202 313636 383610
rect 316024 383202 316084 383610
rect 318472 383202 318532 383610
rect 321056 383202 321116 383610
rect 323368 383202 323428 383610
rect 326088 383610 326170 383670
rect 338438 383670 338498 386275
rect 339726 383670 339786 386275
rect 343794 385308 344414 416898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385308 348134 420618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 385308 351854 388338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 385308 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 350947 385116 351013 385117
rect 350947 385052 350948 385116
rect 351012 385052 351013 385116
rect 350947 385051 351013 385052
rect 350950 383670 351010 385051
rect 338438 383610 338524 383670
rect 326088 383202 326148 383610
rect 338464 383202 338524 383610
rect 339688 383610 339786 383670
rect 350840 383610 351010 383670
rect 339688 383202 339748 383610
rect 350840 383202 350900 383610
rect 220272 381454 220620 381486
rect 220272 381218 220328 381454
rect 220564 381218 220620 381454
rect 220272 381134 220620 381218
rect 220272 380898 220328 381134
rect 220564 380898 220620 381134
rect 220272 380866 220620 380898
rect 356000 381454 356348 381486
rect 356000 381218 356056 381454
rect 356292 381218 356348 381454
rect 356000 381134 356348 381218
rect 356000 380898 356056 381134
rect 356292 380898 356348 381134
rect 356000 380866 356348 380898
rect 220952 363454 221300 363486
rect 220952 363218 221008 363454
rect 221244 363218 221300 363454
rect 220952 363134 221300 363218
rect 220952 362898 221008 363134
rect 221244 362898 221300 363134
rect 220952 362866 221300 362898
rect 355320 363454 355668 363486
rect 355320 363218 355376 363454
rect 355612 363218 355668 363454
rect 355320 363134 355668 363218
rect 355320 362898 355376 363134
rect 355612 362898 355668 363134
rect 355320 362866 355668 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 217547 332756 217613 332757
rect 217547 332692 217548 332756
rect 217612 332692 217613 332756
rect 217547 332691 217613 332692
rect 217363 330988 217429 330989
rect 217363 330924 217364 330988
rect 217428 330924 217429 330988
rect 217363 330923 217429 330924
rect 217179 328132 217245 328133
rect 217179 328068 217180 328132
rect 217244 328068 217245 328132
rect 217179 328067 217245 328068
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 232000 211574 248058
rect 144928 219454 145248 219486
rect 144928 219218 144970 219454
rect 145206 219218 145248 219454
rect 144928 219134 145248 219218
rect 144928 218898 144970 219134
rect 145206 218898 145248 219134
rect 144928 218866 145248 218898
rect 175648 219454 175968 219486
rect 175648 219218 175690 219454
rect 175926 219218 175968 219454
rect 175648 219134 175968 219218
rect 175648 218898 175690 219134
rect 175926 218898 175968 219134
rect 175648 218866 175968 218898
rect 206368 219454 206688 219486
rect 206368 219218 206410 219454
rect 206646 219218 206688 219454
rect 206368 219134 206688 219218
rect 206368 218898 206410 219134
rect 206646 218898 206688 219134
rect 206368 218866 206688 218898
rect 160288 201454 160608 201486
rect 160288 201218 160330 201454
rect 160566 201218 160608 201454
rect 160288 201134 160608 201218
rect 160288 200898 160330 201134
rect 160566 200898 160608 201134
rect 160288 200866 160608 200898
rect 191008 201454 191328 201486
rect 191008 201218 191050 201454
rect 191286 201218 191328 201454
rect 191008 201134 191328 201218
rect 191008 200898 191050 201134
rect 191286 200898 191328 201134
rect 191008 200866 191328 200898
rect 144928 183454 145248 183486
rect 144928 183218 144970 183454
rect 145206 183218 145248 183454
rect 144928 183134 145248 183218
rect 144928 182898 144970 183134
rect 145206 182898 145248 183134
rect 144928 182866 145248 182898
rect 175648 183454 175968 183486
rect 175648 183218 175690 183454
rect 175926 183218 175968 183454
rect 175648 183134 175968 183218
rect 175648 182898 175690 183134
rect 175926 182898 175968 183134
rect 175648 182866 175968 182898
rect 206368 183454 206688 183486
rect 206368 183218 206410 183454
rect 206646 183218 206688 183454
rect 206368 183134 206688 183218
rect 206368 182898 206410 183134
rect 206646 182898 206688 183134
rect 206368 182866 206688 182898
rect 160288 165454 160608 165486
rect 160288 165218 160330 165454
rect 160566 165218 160608 165454
rect 160288 165134 160608 165218
rect 160288 164898 160330 165134
rect 160566 164898 160608 165134
rect 160288 164866 160608 164898
rect 191008 165454 191328 165486
rect 191008 165218 191050 165454
rect 191286 165218 191328 165454
rect 191008 165134 191328 165218
rect 191008 164898 191050 165134
rect 191286 164898 191328 165134
rect 191008 164866 191328 164898
rect 217182 160445 217242 328067
rect 217179 160444 217245 160445
rect 217179 160380 217180 160444
rect 217244 160380 217245 160444
rect 217179 160379 217245 160380
rect 217366 158133 217426 330923
rect 217550 158269 217610 332691
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 236056 299570 236116 300106
rect 237144 299570 237204 300106
rect 238232 299570 238292 300106
rect 239592 299570 239652 300106
rect 236056 299510 236562 299570
rect 217794 291454 218414 298000
rect 219203 297804 219269 297805
rect 219203 297740 219204 297804
rect 219268 297740 219269 297804
rect 219203 297739 219269 297740
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 232000 218414 254898
rect 219206 160445 219266 297739
rect 221514 295174 222134 298000
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 232000 222134 258618
rect 225234 262894 225854 298000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 232000 225854 262338
rect 228954 266614 229574 298000
rect 232451 297668 232517 297669
rect 232451 297604 232452 297668
rect 232516 297604 232517 297668
rect 232451 297603 232517 297604
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 232000 229574 266058
rect 221728 201454 222048 201486
rect 221728 201218 221770 201454
rect 222006 201218 222048 201454
rect 221728 201134 222048 201218
rect 221728 200898 221770 201134
rect 222006 200898 222048 201134
rect 221728 200866 222048 200898
rect 221728 165454 222048 165486
rect 221728 165218 221770 165454
rect 222006 165218 222048 165454
rect 221728 165134 222048 165218
rect 221728 164898 221770 165134
rect 222006 164898 222048 165134
rect 221728 164866 222048 164898
rect 219203 160444 219269 160445
rect 219203 160380 219204 160444
rect 219268 160380 219269 160444
rect 219203 160379 219269 160380
rect 232454 158269 232514 297603
rect 235794 273454 236414 298000
rect 236502 297941 236562 299510
rect 237054 299510 237204 299570
rect 238158 299510 238292 299570
rect 239446 299510 239652 299570
rect 240544 299570 240604 300106
rect 241768 299570 241828 300106
rect 243128 299570 243188 300106
rect 240544 299510 240610 299570
rect 241768 299510 241898 299570
rect 237054 298077 237114 299510
rect 238158 298077 238218 299510
rect 239446 299490 239506 299510
rect 238526 299430 239506 299490
rect 237051 298076 237117 298077
rect 237051 298012 237052 298076
rect 237116 298012 237117 298076
rect 237051 298011 237117 298012
rect 238155 298076 238221 298077
rect 238155 298012 238156 298076
rect 238220 298012 238221 298076
rect 238155 298011 238221 298012
rect 236499 297940 236565 297941
rect 236499 297876 236500 297940
rect 236564 297876 236565 297940
rect 236499 297875 236565 297876
rect 238526 296850 238586 299430
rect 238707 296852 238773 296853
rect 238707 296850 238708 296852
rect 238526 296790 238708 296850
rect 238707 296788 238708 296790
rect 238772 296788 238773 296852
rect 238707 296787 238773 296788
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 232000 236414 236898
rect 239514 277174 240134 298000
rect 240550 297805 240610 299510
rect 241838 298077 241898 299510
rect 242942 299510 243188 299570
rect 244216 299570 244276 300106
rect 245440 299570 245500 300106
rect 246528 299570 246588 300106
rect 244216 299510 244290 299570
rect 245440 299510 245578 299570
rect 241835 298076 241901 298077
rect 241835 298012 241836 298076
rect 241900 298012 241901 298076
rect 241835 298011 241901 298012
rect 240547 297804 240613 297805
rect 240547 297740 240548 297804
rect 240612 297740 240613 297804
rect 240547 297739 240613 297740
rect 242942 297669 243002 299510
rect 242939 297668 243005 297669
rect 242939 297604 242940 297668
rect 243004 297604 243005 297668
rect 242939 297603 243005 297604
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 232000 240134 240618
rect 243234 280894 243854 298000
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 232000 243854 244338
rect 237088 219454 237408 219486
rect 237088 219218 237130 219454
rect 237366 219218 237408 219454
rect 237088 219134 237408 219218
rect 237088 218898 237130 219134
rect 237366 218898 237408 219134
rect 237088 218866 237408 218898
rect 237088 183454 237408 183486
rect 237088 183218 237130 183454
rect 237366 183218 237408 183454
rect 237088 183134 237408 183218
rect 237088 182898 237130 183134
rect 237366 182898 237408 183134
rect 237088 182866 237408 182898
rect 244230 158541 244290 299510
rect 245518 297805 245578 299510
rect 246438 299510 246588 299570
rect 247616 299570 247676 300106
rect 248296 299570 248356 300106
rect 248704 299570 248764 300106
rect 247616 299510 247786 299570
rect 245515 297804 245581 297805
rect 245515 297740 245516 297804
rect 245580 297740 245581 297804
rect 245515 297739 245581 297740
rect 246438 296730 246498 299510
rect 247726 298077 247786 299510
rect 248278 299510 248356 299570
rect 248646 299510 248764 299570
rect 250064 299570 250124 300106
rect 250744 299842 250804 300106
rect 251288 299842 251348 300106
rect 250744 299782 250914 299842
rect 250064 299510 250178 299570
rect 247723 298076 247789 298077
rect 247723 298012 247724 298076
rect 247788 298012 247789 298076
rect 247723 298011 247789 298012
rect 245702 296670 246498 296730
rect 244227 158540 244293 158541
rect 244227 158476 244228 158540
rect 244292 158476 244293 158540
rect 244227 158475 244293 158476
rect 245702 158405 245762 296670
rect 246954 284614 247574 298000
rect 248278 297941 248338 299510
rect 248646 298077 248706 299510
rect 250118 298077 250178 299510
rect 250854 298077 250914 299782
rect 251222 299782 251348 299842
rect 251222 298077 251282 299782
rect 252376 299570 252436 300106
rect 253464 299570 253524 300106
rect 252326 299510 252436 299570
rect 253430 299510 253524 299570
rect 253600 299570 253660 300106
rect 254552 299570 254612 300106
rect 255912 299570 255972 300106
rect 253600 299510 253674 299570
rect 252326 298077 252386 299510
rect 248643 298076 248709 298077
rect 248643 298012 248644 298076
rect 248708 298012 248709 298076
rect 248643 298011 248709 298012
rect 250115 298076 250181 298077
rect 250115 298012 250116 298076
rect 250180 298012 250181 298076
rect 250115 298011 250181 298012
rect 250851 298076 250917 298077
rect 250851 298012 250852 298076
rect 250916 298012 250917 298076
rect 250851 298011 250917 298012
rect 251219 298076 251285 298077
rect 251219 298012 251220 298076
rect 251284 298012 251285 298076
rect 251219 298011 251285 298012
rect 252323 298076 252389 298077
rect 252323 298012 252324 298076
rect 252388 298012 252389 298076
rect 252323 298011 252389 298012
rect 248275 297940 248341 297941
rect 248275 297876 248276 297940
rect 248340 297876 248341 297940
rect 248275 297875 248341 297876
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 232000 247574 248058
rect 252448 201454 252768 201486
rect 252448 201218 252490 201454
rect 252726 201218 252768 201454
rect 252448 201134 252768 201218
rect 252448 200898 252490 201134
rect 252726 200898 252768 201134
rect 252448 200866 252768 200898
rect 252448 165454 252768 165486
rect 252448 165218 252490 165454
rect 252726 165218 252768 165454
rect 252448 165134 252768 165218
rect 252448 164898 252490 165134
rect 252726 164898 252768 165134
rect 252448 164866 252768 164898
rect 245699 158404 245765 158405
rect 245699 158340 245700 158404
rect 245764 158340 245765 158404
rect 245699 158339 245765 158340
rect 217547 158268 217613 158269
rect 217547 158204 217548 158268
rect 217612 158204 217613 158268
rect 217547 158203 217613 158204
rect 232451 158268 232517 158269
rect 232451 158204 232452 158268
rect 232516 158204 232517 158268
rect 232451 158203 232517 158204
rect 253430 158133 253490 299510
rect 253614 298077 253674 299510
rect 254534 299510 254612 299570
rect 255822 299510 255972 299570
rect 256048 299570 256108 300106
rect 257000 299570 257060 300106
rect 258088 299570 258148 300106
rect 258496 299570 258556 300106
rect 256048 299510 256250 299570
rect 253611 298076 253677 298077
rect 253611 298012 253612 298076
rect 253676 298012 253677 298076
rect 253611 298011 253677 298012
rect 253794 291454 254414 298000
rect 254534 297125 254594 299510
rect 254531 297124 254597 297125
rect 254531 297060 254532 297124
rect 254596 297060 254597 297124
rect 254531 297059 254597 297060
rect 255822 296853 255882 299510
rect 256190 296989 256250 299510
rect 256926 299510 257060 299570
rect 258030 299510 258148 299570
rect 258398 299510 258556 299570
rect 259448 299570 259508 300106
rect 260672 299570 260732 300106
rect 261080 299570 261140 300106
rect 261760 299570 261820 300106
rect 262848 299570 262908 300106
rect 263528 299570 263588 300106
rect 263936 299570 263996 300106
rect 265296 299570 265356 300106
rect 265976 299570 266036 300106
rect 266384 299570 266444 300106
rect 267608 299570 267668 300106
rect 259448 299510 259562 299570
rect 256187 296988 256253 296989
rect 256187 296924 256188 296988
rect 256252 296924 256253 296988
rect 256187 296923 256253 296924
rect 256926 296853 256986 299510
rect 258030 298213 258090 299510
rect 258027 298212 258093 298213
rect 258027 298148 258028 298212
rect 258092 298148 258093 298212
rect 258027 298147 258093 298148
rect 255819 296852 255885 296853
rect 255819 296788 255820 296852
rect 255884 296788 255885 296852
rect 255819 296787 255885 296788
rect 256923 296852 256989 296853
rect 256923 296788 256924 296852
rect 256988 296788 256989 296852
rect 256923 296787 256989 296788
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 232000 254414 254898
rect 257514 295174 258134 298000
rect 258398 296853 258458 299510
rect 259502 298077 259562 299510
rect 260606 299510 260732 299570
rect 260974 299510 261140 299570
rect 261710 299510 261820 299570
rect 262814 299510 262908 299570
rect 263366 299510 263588 299570
rect 263918 299510 263996 299570
rect 265206 299510 265356 299570
rect 265942 299510 266036 299570
rect 266310 299510 266444 299570
rect 267598 299510 267668 299570
rect 268288 299570 268348 300106
rect 268696 299570 268756 300106
rect 269784 299570 269844 300106
rect 271008 299842 271068 300106
rect 270910 299782 271068 299842
rect 268288 299510 268394 299570
rect 268696 299510 268762 299570
rect 269784 299510 269866 299570
rect 260606 298077 260666 299510
rect 259499 298076 259565 298077
rect 259499 298012 259500 298076
rect 259564 298012 259565 298076
rect 259499 298011 259565 298012
rect 260603 298076 260669 298077
rect 260603 298012 260604 298076
rect 260668 298012 260669 298076
rect 260603 298011 260669 298012
rect 258579 297668 258645 297669
rect 258579 297604 258580 297668
rect 258644 297604 258645 297668
rect 258579 297603 258645 297604
rect 258395 296852 258461 296853
rect 258395 296788 258396 296852
rect 258460 296788 258461 296852
rect 258395 296787 258461 296788
rect 258582 296170 258642 297603
rect 258947 297532 259013 297533
rect 258947 297468 258948 297532
rect 259012 297468 259013 297532
rect 258947 297467 259013 297468
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 232000 258134 258618
rect 258214 296110 258642 296170
rect 258214 171150 258274 296110
rect 258395 296036 258461 296037
rect 258395 295972 258396 296036
rect 258460 295972 258461 296036
rect 258395 295971 258461 295972
rect 258398 180810 258458 295971
rect 258950 294810 259010 297467
rect 259499 297260 259565 297261
rect 259499 297196 259500 297260
rect 259564 297196 259565 297260
rect 259499 297195 259565 297196
rect 259131 297124 259197 297125
rect 259131 297060 259132 297124
rect 259196 297060 259197 297124
rect 259131 297059 259197 297060
rect 258582 294750 259010 294810
rect 258582 190470 258642 294750
rect 259134 292590 259194 297059
rect 258766 292530 259194 292590
rect 258766 209790 258826 292530
rect 258766 209730 259378 209790
rect 259318 197573 259378 209730
rect 259315 197572 259381 197573
rect 259315 197508 259316 197572
rect 259380 197508 259381 197572
rect 259315 197507 259381 197508
rect 258582 190410 259378 190470
rect 259318 186421 259378 190410
rect 259315 186420 259381 186421
rect 259315 186356 259316 186420
rect 259380 186356 259381 186420
rect 259315 186355 259381 186356
rect 258398 180750 259378 180810
rect 259318 175269 259378 180750
rect 259315 175268 259381 175269
rect 259315 175204 259316 175268
rect 259380 175204 259381 175268
rect 259315 175203 259381 175204
rect 258214 171090 259378 171150
rect 259318 164253 259378 171090
rect 259502 170781 259562 297195
rect 260974 296853 261034 299510
rect 261710 298213 261770 299510
rect 261707 298212 261773 298213
rect 261707 298148 261708 298212
rect 261772 298148 261773 298212
rect 261707 298147 261773 298148
rect 260971 296852 261037 296853
rect 260971 296788 260972 296852
rect 261036 296788 261037 296852
rect 260971 296787 261037 296788
rect 261234 262894 261854 298000
rect 262814 296853 262874 299510
rect 263366 298074 263426 299510
rect 263547 298076 263613 298077
rect 263547 298074 263548 298076
rect 263366 298014 263548 298074
rect 263547 298012 263548 298014
rect 263612 298012 263613 298076
rect 263547 298011 263613 298012
rect 263918 297941 263978 299510
rect 265206 298213 265266 299510
rect 265203 298212 265269 298213
rect 265203 298148 265204 298212
rect 265268 298148 265269 298212
rect 265203 298147 265269 298148
rect 265942 298077 266002 299510
rect 266310 298077 266370 299510
rect 265939 298076 266005 298077
rect 265939 298012 265940 298076
rect 266004 298012 266005 298076
rect 265939 298011 266005 298012
rect 266307 298076 266373 298077
rect 266307 298012 266308 298076
rect 266372 298012 266373 298076
rect 266307 298011 266373 298012
rect 263915 297940 263981 297941
rect 263915 297876 263916 297940
rect 263980 297876 263981 297940
rect 263915 297875 263981 297876
rect 262811 296852 262877 296853
rect 262811 296788 262812 296852
rect 262876 296788 262877 296852
rect 262811 296787 262877 296788
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 259683 239460 259749 239461
rect 259683 239396 259684 239460
rect 259748 239396 259749 239460
rect 259683 239395 259749 239396
rect 259686 184925 259746 239395
rect 261234 232000 261854 262338
rect 264954 266614 265574 298000
rect 267598 297941 267658 299510
rect 268334 297941 268394 299510
rect 268702 298077 268762 299510
rect 269806 298077 269866 299510
rect 270910 298077 270970 299782
rect 271144 299570 271204 300106
rect 272232 299570 272292 300106
rect 273320 299570 273380 300106
rect 273592 299842 273652 300106
rect 271094 299510 271204 299570
rect 272198 299510 272292 299570
rect 273302 299510 273380 299570
rect 273486 299782 273652 299842
rect 268699 298076 268765 298077
rect 268699 298012 268700 298076
rect 268764 298012 268765 298076
rect 268699 298011 268765 298012
rect 269803 298076 269869 298077
rect 269803 298012 269804 298076
rect 269868 298012 269869 298076
rect 269803 298011 269869 298012
rect 270907 298076 270973 298077
rect 270907 298012 270908 298076
rect 270972 298012 270973 298076
rect 270907 298011 270973 298012
rect 271094 297941 271154 299510
rect 272198 298213 272258 299510
rect 272195 298212 272261 298213
rect 272195 298148 272196 298212
rect 272260 298148 272261 298212
rect 272195 298147 272261 298148
rect 273302 298077 273362 299510
rect 273299 298076 273365 298077
rect 273299 298012 273300 298076
rect 273364 298012 273365 298076
rect 273299 298011 273365 298012
rect 267595 297940 267661 297941
rect 267595 297876 267596 297940
rect 267660 297876 267661 297940
rect 267595 297875 267661 297876
rect 268331 297940 268397 297941
rect 268331 297876 268332 297940
rect 268396 297876 268397 297940
rect 268331 297875 268397 297876
rect 271091 297940 271157 297941
rect 271091 297876 271092 297940
rect 271156 297876 271157 297940
rect 271091 297875 271157 297876
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 262811 230212 262877 230213
rect 262811 230148 262812 230212
rect 262876 230148 262877 230212
rect 262811 230147 262877 230148
rect 262443 230076 262509 230077
rect 262443 230012 262444 230076
rect 262508 230012 262509 230076
rect 262443 230011 262509 230012
rect 262259 229940 262325 229941
rect 262259 229876 262260 229940
rect 262324 229876 262325 229940
rect 262259 229875 262325 229876
rect 259683 184924 259749 184925
rect 259683 184860 259684 184924
rect 259748 184860 259749 184924
rect 259683 184859 259749 184860
rect 259499 170780 259565 170781
rect 259499 170716 259500 170780
rect 259564 170716 259565 170780
rect 259499 170715 259565 170716
rect 262262 167653 262322 229875
rect 262446 177309 262506 230011
rect 262627 229668 262693 229669
rect 262627 229604 262628 229668
rect 262692 229604 262693 229668
rect 262627 229603 262693 229604
rect 262630 183565 262690 229603
rect 262814 194581 262874 230147
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 262811 194580 262877 194581
rect 262811 194516 262812 194580
rect 262876 194516 262877 194580
rect 262811 194515 262877 194516
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 262627 183564 262693 183565
rect 262627 183500 262628 183564
rect 262692 183500 262693 183564
rect 262627 183499 262693 183500
rect 262443 177308 262509 177309
rect 262443 177244 262444 177308
rect 262508 177244 262509 177308
rect 262443 177243 262509 177244
rect 262259 167652 262325 167653
rect 262259 167588 262260 167652
rect 262324 167588 262325 167652
rect 262259 167587 262325 167588
rect 259315 164252 259381 164253
rect 259315 164188 259316 164252
rect 259380 164188 259381 164252
rect 259315 164187 259381 164188
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 217363 158132 217429 158133
rect 217363 158068 217364 158132
rect 217428 158068 217429 158132
rect 217363 158067 217429 158068
rect 253427 158132 253493 158133
rect 253427 158068 253428 158132
rect 253492 158068 253493 158132
rect 253427 158067 253493 158068
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 129963 157996 130029 157997
rect 129963 157932 129964 157996
rect 130028 157932 130029 157996
rect 129963 157931 130029 157932
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 133174 132134 158000
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 136894 135854 158000
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 140614 139574 158000
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 147454 146414 158000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 151174 150134 158000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 154894 153854 158000
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 122614 157574 158000
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 129454 164414 158000
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 133174 168134 158000
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 136894 171854 158000
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 140614 175574 158000
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 147454 182414 158000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 151174 186134 158000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 154894 189854 158000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 122614 193574 158000
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 129454 200414 158000
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 133174 204134 158000
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 136894 207854 158000
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 140614 211574 158000
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 151174 222134 158000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 154894 225854 158000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 122614 229574 158000
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 129454 236414 158000
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 133174 240134 158000
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 136894 243854 158000
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 140614 247574 158000
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 158000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 257514 151174 258134 158000
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 122000 258134 150618
rect 261234 154894 261854 158000
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 122000 261854 154338
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 122000 265574 122058
rect 271794 273454 272414 298000
rect 273486 297941 273546 299782
rect 274408 299570 274468 300106
rect 275768 299842 275828 300106
rect 274406 299510 274468 299570
rect 275694 299782 275828 299842
rect 273483 297940 273549 297941
rect 273483 297876 273484 297940
rect 273548 297876 273549 297940
rect 273483 297875 273549 297876
rect 274406 297805 274466 299510
rect 275694 298213 275754 299782
rect 276040 299570 276100 300106
rect 276992 299570 277052 300106
rect 276040 299510 276122 299570
rect 276062 298213 276122 299510
rect 276982 299510 277052 299570
rect 278080 299570 278140 300106
rect 278488 299570 278548 300106
rect 279168 299570 279228 300106
rect 280936 299570 280996 300106
rect 283520 299570 283580 300106
rect 278080 299510 278146 299570
rect 275691 298212 275757 298213
rect 275691 298148 275692 298212
rect 275756 298148 275757 298212
rect 275691 298147 275757 298148
rect 276059 298212 276125 298213
rect 276059 298148 276060 298212
rect 276124 298148 276125 298212
rect 276059 298147 276125 298148
rect 276982 298077 277042 299510
rect 276979 298076 277045 298077
rect 276979 298012 276980 298076
rect 277044 298012 277045 298076
rect 276979 298011 277045 298012
rect 274403 297804 274469 297805
rect 274403 297740 274404 297804
rect 274468 297740 274469 297804
rect 274403 297739 274469 297740
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 122000 272414 128898
rect 275514 277174 276134 298000
rect 278086 296989 278146 299510
rect 278454 299510 278548 299570
rect 279006 299510 279228 299570
rect 280846 299510 280996 299570
rect 283422 299510 283580 299570
rect 285968 299570 286028 300106
rect 288280 299570 288340 300106
rect 291000 299570 291060 300106
rect 293448 299570 293508 300106
rect 285968 299510 286058 299570
rect 278454 298077 278514 299510
rect 279006 298077 279066 299510
rect 280846 298077 280906 299510
rect 283422 298213 283482 299510
rect 283419 298212 283485 298213
rect 283419 298148 283420 298212
rect 283484 298148 283485 298212
rect 283419 298147 283485 298148
rect 285998 298077 286058 299510
rect 288206 299510 288340 299570
rect 290966 299510 291060 299570
rect 293358 299510 293508 299570
rect 295896 299570 295956 300106
rect 298480 299570 298540 300106
rect 300928 299570 300988 300106
rect 303512 299570 303572 300106
rect 305960 299570 306020 300106
rect 295896 299510 295994 299570
rect 298480 299510 298570 299570
rect 288206 298077 288266 299510
rect 290966 298077 291026 299510
rect 293358 298077 293418 299510
rect 295934 298077 295994 299510
rect 298510 298077 298570 299510
rect 300902 299510 300988 299570
rect 303478 299510 303572 299570
rect 305870 299510 306020 299570
rect 308544 299570 308604 300106
rect 310992 299570 311052 300106
rect 313440 299570 313500 300106
rect 315888 299570 315948 300106
rect 318472 299570 318532 300106
rect 308544 299510 308690 299570
rect 310992 299510 311082 299570
rect 300902 298213 300962 299510
rect 300899 298212 300965 298213
rect 300899 298148 300900 298212
rect 300964 298148 300965 298212
rect 300899 298147 300965 298148
rect 303478 298077 303538 299510
rect 305870 298077 305930 299510
rect 308630 298077 308690 299510
rect 311022 298077 311082 299510
rect 313414 299510 313500 299570
rect 315806 299510 315948 299570
rect 318382 299510 318532 299570
rect 320920 299570 320980 300106
rect 323368 299570 323428 300106
rect 325952 299570 326012 300106
rect 343224 299570 343284 300106
rect 320920 299510 321018 299570
rect 313414 298077 313474 299510
rect 315806 298213 315866 299510
rect 315803 298212 315869 298213
rect 315803 298148 315804 298212
rect 315868 298148 315869 298212
rect 315803 298147 315869 298148
rect 318382 298077 318442 299510
rect 320958 298077 321018 299510
rect 323350 299510 323428 299570
rect 325926 299510 326012 299570
rect 343222 299510 343284 299570
rect 343360 299570 343420 300106
rect 343360 299510 343466 299570
rect 323350 298077 323410 299510
rect 325926 298213 325986 299510
rect 325923 298212 325989 298213
rect 325923 298148 325924 298212
rect 325988 298148 325989 298212
rect 325923 298147 325989 298148
rect 343222 298077 343282 299510
rect 343406 298077 343466 299510
rect 278451 298076 278517 298077
rect 278451 298012 278452 298076
rect 278516 298012 278517 298076
rect 278451 298011 278517 298012
rect 279003 298076 279069 298077
rect 279003 298012 279004 298076
rect 279068 298012 279069 298076
rect 279003 298011 279069 298012
rect 280843 298076 280909 298077
rect 280843 298012 280844 298076
rect 280908 298012 280909 298076
rect 280843 298011 280909 298012
rect 285995 298076 286061 298077
rect 285995 298012 285996 298076
rect 286060 298012 286061 298076
rect 285995 298011 286061 298012
rect 288203 298076 288269 298077
rect 288203 298012 288204 298076
rect 288268 298012 288269 298076
rect 288203 298011 288269 298012
rect 290963 298076 291029 298077
rect 290963 298012 290964 298076
rect 291028 298012 291029 298076
rect 290963 298011 291029 298012
rect 293355 298076 293421 298077
rect 293355 298012 293356 298076
rect 293420 298012 293421 298076
rect 293355 298011 293421 298012
rect 295931 298076 295997 298077
rect 295931 298012 295932 298076
rect 295996 298012 295997 298076
rect 295931 298011 295997 298012
rect 298507 298076 298573 298077
rect 298507 298012 298508 298076
rect 298572 298012 298573 298076
rect 298507 298011 298573 298012
rect 303475 298076 303541 298077
rect 303475 298012 303476 298076
rect 303540 298012 303541 298076
rect 303475 298011 303541 298012
rect 305867 298076 305933 298077
rect 305867 298012 305868 298076
rect 305932 298012 305933 298076
rect 305867 298011 305933 298012
rect 308627 298076 308693 298077
rect 308627 298012 308628 298076
rect 308692 298012 308693 298076
rect 308627 298011 308693 298012
rect 311019 298076 311085 298077
rect 311019 298012 311020 298076
rect 311084 298012 311085 298076
rect 311019 298011 311085 298012
rect 313411 298076 313477 298077
rect 313411 298012 313412 298076
rect 313476 298012 313477 298076
rect 313411 298011 313477 298012
rect 318379 298076 318445 298077
rect 318379 298012 318380 298076
rect 318444 298012 318445 298076
rect 318379 298011 318445 298012
rect 320955 298076 321021 298077
rect 320955 298012 320956 298076
rect 321020 298012 321021 298076
rect 320955 298011 321021 298012
rect 323347 298076 323413 298077
rect 323347 298012 323348 298076
rect 323412 298012 323413 298076
rect 323347 298011 323413 298012
rect 343219 298076 343285 298077
rect 343219 298012 343220 298076
rect 343284 298012 343285 298076
rect 343219 298011 343285 298012
rect 343403 298076 343469 298077
rect 343403 298012 343404 298076
rect 343468 298012 343469 298076
rect 343403 298011 343469 298012
rect 278083 296988 278149 296989
rect 278083 296924 278084 296988
rect 278148 296924 278149 296988
rect 278083 296923 278149 296924
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 122000 276134 132618
rect 279234 280894 279854 298000
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 122000 279854 136338
rect 282954 284614 283574 298000
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 122000 283574 140058
rect 289794 291454 290414 298000
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 122000 290414 146898
rect 293514 295174 294134 298000
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 122000 294134 150618
rect 297234 262894 297854 298000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 122000 297854 154338
rect 300954 266614 301574 298000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 122000 301574 122058
rect 307794 273454 308414 298000
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 122000 308414 128898
rect 311514 277174 312134 298000
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 122000 312134 132618
rect 315234 280894 315854 298000
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 122000 315854 136338
rect 318954 284614 319574 298000
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 122000 319574 140058
rect 325794 291454 326414 298000
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 122000 326414 146898
rect 329514 295174 330134 298000
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 122000 330134 150618
rect 333234 262894 333854 298000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 122000 333854 154338
rect 336954 266614 337574 298000
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 122000 337574 122058
rect 343794 273454 344414 298000
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 264208 111454 264528 111486
rect 264208 111218 264250 111454
rect 264486 111218 264528 111454
rect 264208 111134 264528 111218
rect 264208 110898 264250 111134
rect 264486 110898 264528 111134
rect 264208 110866 264528 110898
rect 294928 111454 295248 111486
rect 294928 111218 294970 111454
rect 295206 111218 295248 111454
rect 294928 111134 295248 111218
rect 294928 110898 294970 111134
rect 295206 110898 295248 111134
rect 294928 110866 295248 110898
rect 325648 111454 325968 111486
rect 325648 111218 325690 111454
rect 325926 111218 325968 111454
rect 325648 111134 325968 111218
rect 325648 110898 325690 111134
rect 325926 110898 325968 111134
rect 325648 110866 325968 110898
rect 279568 93454 279888 93486
rect 279568 93218 279610 93454
rect 279846 93218 279888 93454
rect 279568 93134 279888 93218
rect 279568 92898 279610 93134
rect 279846 92898 279888 93134
rect 279568 92866 279888 92898
rect 310288 93454 310608 93486
rect 310288 93218 310330 93454
rect 310566 93218 310608 93454
rect 310288 93134 310608 93218
rect 310288 92898 310330 93134
rect 310566 92898 310608 93134
rect 310288 92866 310608 92898
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 264208 75454 264528 75486
rect 264208 75218 264250 75454
rect 264486 75218 264528 75454
rect 264208 75134 264528 75218
rect 264208 74898 264250 75134
rect 264486 74898 264528 75134
rect 264208 74866 264528 74898
rect 294928 75454 295248 75486
rect 294928 75218 294970 75454
rect 295206 75218 295248 75454
rect 294928 75134 295248 75218
rect 294928 74898 294970 75134
rect 295206 74898 295248 75134
rect 294928 74866 295248 74898
rect 325648 75454 325968 75486
rect 325648 75218 325690 75454
rect 325926 75218 325968 75454
rect 325648 75134 325968 75218
rect 325648 74898 325690 75134
rect 325926 74898 325968 75134
rect 325648 74866 325968 74898
rect 279568 57454 279888 57486
rect 279568 57218 279610 57454
rect 279846 57218 279888 57454
rect 279568 57134 279888 57218
rect 279568 56898 279610 57134
rect 279846 56898 279888 57134
rect 279568 56866 279888 56898
rect 310288 57454 310608 57486
rect 310288 57218 310330 57454
rect 310566 57218 310608 57454
rect 310288 57134 310608 57218
rect 310288 56898 310330 57134
rect 310566 56898 310608 57134
rect 310288 56866 310608 56898
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 38000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 38000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 38000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 38000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 38000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 38000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 38000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 3454 290414 38000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 38000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 38000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 38000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 38000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 38000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 38000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 38000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 3454 326414 38000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 38000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 38000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 38000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 277174 348134 298000
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 280894 351854 298000
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 284614 355574 298000
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 552000 380414 560898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 552000 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 552000 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 552000 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 552000 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 552000 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 552000 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 552000 409574 554058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 552000 416414 560898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 552000 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 552000 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 552000 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 552000 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 552000 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 552000 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 552000 445574 554058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 552000 452414 560898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 552000 456134 564618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 552000 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 552000 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 552000 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 552000 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 552000 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 552000 481574 554058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 552000 488414 560898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 552000 492134 564618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 552000 495854 568338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 552000 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 552000 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 552000 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 552000 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 552000 517574 554058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 552000 524414 560898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 552000 528134 564618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 552000 531854 568338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 384208 543454 384528 543486
rect 384208 543218 384250 543454
rect 384486 543218 384528 543454
rect 384208 543134 384528 543218
rect 384208 542898 384250 543134
rect 384486 542898 384528 543134
rect 384208 542866 384528 542898
rect 414928 543454 415248 543486
rect 414928 543218 414970 543454
rect 415206 543218 415248 543454
rect 414928 543134 415248 543218
rect 414928 542898 414970 543134
rect 415206 542898 415248 543134
rect 414928 542866 415248 542898
rect 445648 543454 445968 543486
rect 445648 543218 445690 543454
rect 445926 543218 445968 543454
rect 445648 543134 445968 543218
rect 445648 542898 445690 543134
rect 445926 542898 445968 543134
rect 445648 542866 445968 542898
rect 476368 543454 476688 543486
rect 476368 543218 476410 543454
rect 476646 543218 476688 543454
rect 476368 543134 476688 543218
rect 476368 542898 476410 543134
rect 476646 542898 476688 543134
rect 476368 542866 476688 542898
rect 507088 543454 507408 543486
rect 507088 543218 507130 543454
rect 507366 543218 507408 543454
rect 507088 543134 507408 543218
rect 507088 542898 507130 543134
rect 507366 542898 507408 543134
rect 507088 542866 507408 542898
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 399568 525454 399888 525486
rect 399568 525218 399610 525454
rect 399846 525218 399888 525454
rect 399568 525134 399888 525218
rect 399568 524898 399610 525134
rect 399846 524898 399888 525134
rect 399568 524866 399888 524898
rect 430288 525454 430608 525486
rect 430288 525218 430330 525454
rect 430566 525218 430608 525454
rect 430288 525134 430608 525218
rect 430288 524898 430330 525134
rect 430566 524898 430608 525134
rect 430288 524866 430608 524898
rect 461008 525454 461328 525486
rect 461008 525218 461050 525454
rect 461286 525218 461328 525454
rect 461008 525134 461328 525218
rect 461008 524898 461050 525134
rect 461286 524898 461328 525134
rect 461008 524866 461328 524898
rect 491728 525454 492048 525486
rect 491728 525218 491770 525454
rect 492006 525218 492048 525454
rect 491728 525134 492048 525218
rect 491728 524898 491770 525134
rect 492006 524898 492048 525134
rect 491728 524866 492048 524898
rect 522448 525454 522768 525486
rect 522448 525218 522490 525454
rect 522726 525218 522768 525454
rect 522448 525134 522768 525218
rect 522448 524898 522490 525134
rect 522726 524898 522768 525134
rect 522448 524866 522768 524898
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 384208 507454 384528 507486
rect 384208 507218 384250 507454
rect 384486 507218 384528 507454
rect 384208 507134 384528 507218
rect 384208 506898 384250 507134
rect 384486 506898 384528 507134
rect 384208 506866 384528 506898
rect 414928 507454 415248 507486
rect 414928 507218 414970 507454
rect 415206 507218 415248 507454
rect 414928 507134 415248 507218
rect 414928 506898 414970 507134
rect 415206 506898 415248 507134
rect 414928 506866 415248 506898
rect 445648 507454 445968 507486
rect 445648 507218 445690 507454
rect 445926 507218 445968 507454
rect 445648 507134 445968 507218
rect 445648 506898 445690 507134
rect 445926 506898 445968 507134
rect 445648 506866 445968 506898
rect 476368 507454 476688 507486
rect 476368 507218 476410 507454
rect 476646 507218 476688 507454
rect 476368 507134 476688 507218
rect 476368 506898 476410 507134
rect 476646 506898 476688 507134
rect 476368 506866 476688 506898
rect 507088 507454 507408 507486
rect 507088 507218 507130 507454
rect 507366 507218 507408 507454
rect 507088 507134 507408 507218
rect 507088 506898 507130 507134
rect 507366 506898 507408 507134
rect 507088 506866 507408 506898
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 399568 489454 399888 489486
rect 399568 489218 399610 489454
rect 399846 489218 399888 489454
rect 399568 489134 399888 489218
rect 399568 488898 399610 489134
rect 399846 488898 399888 489134
rect 399568 488866 399888 488898
rect 430288 489454 430608 489486
rect 430288 489218 430330 489454
rect 430566 489218 430608 489454
rect 430288 489134 430608 489218
rect 430288 488898 430330 489134
rect 430566 488898 430608 489134
rect 430288 488866 430608 488898
rect 461008 489454 461328 489486
rect 461008 489218 461050 489454
rect 461286 489218 461328 489454
rect 461008 489134 461328 489218
rect 461008 488898 461050 489134
rect 461286 488898 461328 489134
rect 461008 488866 461328 488898
rect 491728 489454 492048 489486
rect 491728 489218 491770 489454
rect 492006 489218 492048 489454
rect 491728 489134 492048 489218
rect 491728 488898 491770 489134
rect 492006 488898 492048 489134
rect 491728 488866 492048 488898
rect 522448 489454 522768 489486
rect 522448 489218 522490 489454
rect 522726 489218 522768 489454
rect 522448 489134 522768 489218
rect 522448 488898 522490 489134
rect 522726 488898 522768 489134
rect 522448 488866 522768 488898
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 384208 471454 384528 471486
rect 384208 471218 384250 471454
rect 384486 471218 384528 471454
rect 384208 471134 384528 471218
rect 384208 470898 384250 471134
rect 384486 470898 384528 471134
rect 384208 470866 384528 470898
rect 414928 471454 415248 471486
rect 414928 471218 414970 471454
rect 415206 471218 415248 471454
rect 414928 471134 415248 471218
rect 414928 470898 414970 471134
rect 415206 470898 415248 471134
rect 414928 470866 415248 470898
rect 445648 471454 445968 471486
rect 445648 471218 445690 471454
rect 445926 471218 445968 471454
rect 445648 471134 445968 471218
rect 445648 470898 445690 471134
rect 445926 470898 445968 471134
rect 445648 470866 445968 470898
rect 476368 471454 476688 471486
rect 476368 471218 476410 471454
rect 476646 471218 476688 471454
rect 476368 471134 476688 471218
rect 476368 470898 476410 471134
rect 476646 470898 476688 471134
rect 476368 470866 476688 470898
rect 507088 471454 507408 471486
rect 507088 471218 507130 471454
rect 507366 471218 507408 471454
rect 507088 471134 507408 471218
rect 507088 470898 507130 471134
rect 507366 470898 507408 471134
rect 507088 470866 507408 470898
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 399568 453454 399888 453486
rect 399568 453218 399610 453454
rect 399846 453218 399888 453454
rect 399568 453134 399888 453218
rect 399568 452898 399610 453134
rect 399846 452898 399888 453134
rect 399568 452866 399888 452898
rect 430288 453454 430608 453486
rect 430288 453218 430330 453454
rect 430566 453218 430608 453454
rect 430288 453134 430608 453218
rect 430288 452898 430330 453134
rect 430566 452898 430608 453134
rect 430288 452866 430608 452898
rect 461008 453454 461328 453486
rect 461008 453218 461050 453454
rect 461286 453218 461328 453454
rect 461008 453134 461328 453218
rect 461008 452898 461050 453134
rect 461286 452898 461328 453134
rect 461008 452866 461328 452898
rect 491728 453454 492048 453486
rect 491728 453218 491770 453454
rect 492006 453218 492048 453454
rect 491728 453134 492048 453218
rect 491728 452898 491770 453134
rect 492006 452898 492048 453134
rect 491728 452866 492048 452898
rect 522448 453454 522768 453486
rect 522448 453218 522490 453454
rect 522726 453218 522768 453454
rect 522448 453134 522768 453218
rect 522448 452898 522490 453134
rect 522726 452898 522768 453134
rect 522448 452866 522768 452898
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 417454 380414 438000
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 421174 384134 438000
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 424894 387854 438000
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 428614 391574 438000
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 435454 398414 438000
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 403174 402134 438000
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 406894 405854 438000
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 410614 409574 438000
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 417454 416414 438000
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 421174 420134 438000
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 424894 423854 438000
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 428614 427574 438000
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 435454 434414 438000
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 403174 438134 438000
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 406894 441854 438000
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 410614 445574 438000
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 417454 452414 438000
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 421174 456134 438000
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 424894 459854 438000
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 428614 463574 438000
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 435454 470414 438000
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 403174 474134 438000
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 406894 477854 438000
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 410614 481574 438000
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 417454 488414 438000
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 421174 492134 438000
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 424894 495854 438000
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 428614 499574 438000
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 435454 506414 438000
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 403174 510134 438000
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 406894 513854 438000
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 410614 517574 438000
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 417454 524414 438000
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 421174 528134 438000
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 424894 531854 438000
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 149610 489218 149846 489454
rect 149610 488898 149846 489134
rect 180330 489218 180566 489454
rect 180330 488898 180566 489134
rect 211050 489218 211286 489454
rect 211050 488898 211286 489134
rect 241770 489218 242006 489454
rect 241770 488898 242006 489134
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 134250 471218 134486 471454
rect 134250 470898 134486 471134
rect 164970 471218 165206 471454
rect 164970 470898 165206 471134
rect 195690 471218 195926 471454
rect 195690 470898 195926 471134
rect 226410 471218 226646 471454
rect 226410 470898 226646 471134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 40328 381218 40564 381454
rect 40328 380898 40564 381134
rect 176056 381218 176292 381454
rect 176056 380898 176292 381134
rect 41008 363218 41244 363454
rect 41008 362898 41244 363134
rect 175376 363218 175612 363454
rect 175376 362898 175612 363134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 40328 345218 40564 345454
rect 40328 344898 40564 345134
rect 176056 345218 176292 345454
rect 176056 344898 176292 345134
rect 41008 327218 41244 327454
rect 41008 326898 41244 327134
rect 175376 327218 175612 327454
rect 175376 326898 175612 327134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 40328 309218 40564 309454
rect 40328 308898 40564 309134
rect 176056 309218 176292 309454
rect 176056 308898 176292 309134
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 114250 219218 114486 219454
rect 114250 218898 114486 219134
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 129610 201218 129846 201454
rect 129610 200898 129846 201134
rect 114250 183218 114486 183454
rect 114250 182898 114486 183134
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 129610 165218 129846 165454
rect 129610 164898 129846 165134
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 220328 381218 220564 381454
rect 220328 380898 220564 381134
rect 356056 381218 356292 381454
rect 356056 380898 356292 381134
rect 221008 363218 221244 363454
rect 221008 362898 221244 363134
rect 355376 363218 355612 363454
rect 355376 362898 355612 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 144970 219218 145206 219454
rect 144970 218898 145206 219134
rect 175690 219218 175926 219454
rect 175690 218898 175926 219134
rect 206410 219218 206646 219454
rect 206410 218898 206646 219134
rect 160330 201218 160566 201454
rect 160330 200898 160566 201134
rect 191050 201218 191286 201454
rect 191050 200898 191286 201134
rect 144970 183218 145206 183454
rect 144970 182898 145206 183134
rect 175690 183218 175926 183454
rect 175690 182898 175926 183134
rect 206410 183218 206646 183454
rect 206410 182898 206646 183134
rect 160330 165218 160566 165454
rect 160330 164898 160566 165134
rect 191050 165218 191286 165454
rect 191050 164898 191286 165134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 221770 201218 222006 201454
rect 221770 200898 222006 201134
rect 221770 165218 222006 165454
rect 221770 164898 222006 165134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 237130 219218 237366 219454
rect 237130 218898 237366 219134
rect 237130 183218 237366 183454
rect 237130 182898 237366 183134
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 252490 201218 252726 201454
rect 252490 200898 252726 201134
rect 252490 165218 252726 165454
rect 252490 164898 252726 165134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 264250 111218 264486 111454
rect 264250 110898 264486 111134
rect 294970 111218 295206 111454
rect 294970 110898 295206 111134
rect 325690 111218 325926 111454
rect 325690 110898 325926 111134
rect 279610 93218 279846 93454
rect 279610 92898 279846 93134
rect 310330 93218 310566 93454
rect 310330 92898 310566 93134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 264250 75218 264486 75454
rect 264250 74898 264486 75134
rect 294970 75218 295206 75454
rect 294970 74898 295206 75134
rect 325690 75218 325926 75454
rect 325690 74898 325926 75134
rect 279610 57218 279846 57454
rect 279610 56898 279846 57134
rect 310330 57218 310566 57454
rect 310330 56898 310566 57134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 384250 543218 384486 543454
rect 384250 542898 384486 543134
rect 414970 543218 415206 543454
rect 414970 542898 415206 543134
rect 445690 543218 445926 543454
rect 445690 542898 445926 543134
rect 476410 543218 476646 543454
rect 476410 542898 476646 543134
rect 507130 543218 507366 543454
rect 507130 542898 507366 543134
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 399610 525218 399846 525454
rect 399610 524898 399846 525134
rect 430330 525218 430566 525454
rect 430330 524898 430566 525134
rect 461050 525218 461286 525454
rect 461050 524898 461286 525134
rect 491770 525218 492006 525454
rect 491770 524898 492006 525134
rect 522490 525218 522726 525454
rect 522490 524898 522726 525134
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 384250 507218 384486 507454
rect 384250 506898 384486 507134
rect 414970 507218 415206 507454
rect 414970 506898 415206 507134
rect 445690 507218 445926 507454
rect 445690 506898 445926 507134
rect 476410 507218 476646 507454
rect 476410 506898 476646 507134
rect 507130 507218 507366 507454
rect 507130 506898 507366 507134
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 399610 489218 399846 489454
rect 399610 488898 399846 489134
rect 430330 489218 430566 489454
rect 430330 488898 430566 489134
rect 461050 489218 461286 489454
rect 461050 488898 461286 489134
rect 491770 489218 492006 489454
rect 491770 488898 492006 489134
rect 522490 489218 522726 489454
rect 522490 488898 522726 489134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 384250 471218 384486 471454
rect 384250 470898 384486 471134
rect 414970 471218 415206 471454
rect 414970 470898 415206 471134
rect 445690 471218 445926 471454
rect 445690 470898 445926 471134
rect 476410 471218 476646 471454
rect 476410 470898 476646 471134
rect 507130 471218 507366 471454
rect 507130 470898 507366 471134
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 399610 453218 399846 453454
rect 399610 452898 399846 453134
rect 430330 453218 430566 453454
rect 430330 452898 430566 453134
rect 461050 453218 461286 453454
rect 461050 452898 461286 453134
rect 491770 453218 492006 453454
rect 491770 452898 492006 453134
rect 522490 453218 522726 453454
rect 522490 452898 522726 453134
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 384250 543454
rect 384486 543218 414970 543454
rect 415206 543218 445690 543454
rect 445926 543218 476410 543454
rect 476646 543218 507130 543454
rect 507366 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 384250 543134
rect 384486 542898 414970 543134
rect 415206 542898 445690 543134
rect 445926 542898 476410 543134
rect 476646 542898 507130 543134
rect 507366 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 399610 525454
rect 399846 525218 430330 525454
rect 430566 525218 461050 525454
rect 461286 525218 491770 525454
rect 492006 525218 522490 525454
rect 522726 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 399610 525134
rect 399846 524898 430330 525134
rect 430566 524898 461050 525134
rect 461286 524898 491770 525134
rect 492006 524898 522490 525134
rect 522726 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 384250 507454
rect 384486 507218 414970 507454
rect 415206 507218 445690 507454
rect 445926 507218 476410 507454
rect 476646 507218 507130 507454
rect 507366 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 384250 507134
rect 384486 506898 414970 507134
rect 415206 506898 445690 507134
rect 445926 506898 476410 507134
rect 476646 506898 507130 507134
rect 507366 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 149610 489454
rect 149846 489218 180330 489454
rect 180566 489218 211050 489454
rect 211286 489218 241770 489454
rect 242006 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 399610 489454
rect 399846 489218 430330 489454
rect 430566 489218 461050 489454
rect 461286 489218 491770 489454
rect 492006 489218 522490 489454
rect 522726 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 149610 489134
rect 149846 488898 180330 489134
rect 180566 488898 211050 489134
rect 211286 488898 241770 489134
rect 242006 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 399610 489134
rect 399846 488898 430330 489134
rect 430566 488898 461050 489134
rect 461286 488898 491770 489134
rect 492006 488898 522490 489134
rect 522726 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 134250 471454
rect 134486 471218 164970 471454
rect 165206 471218 195690 471454
rect 195926 471218 226410 471454
rect 226646 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 384250 471454
rect 384486 471218 414970 471454
rect 415206 471218 445690 471454
rect 445926 471218 476410 471454
rect 476646 471218 507130 471454
rect 507366 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 134250 471134
rect 134486 470898 164970 471134
rect 165206 470898 195690 471134
rect 195926 470898 226410 471134
rect 226646 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 384250 471134
rect 384486 470898 414970 471134
rect 415206 470898 445690 471134
rect 445926 470898 476410 471134
rect 476646 470898 507130 471134
rect 507366 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 399610 453454
rect 399846 453218 430330 453454
rect 430566 453218 461050 453454
rect 461286 453218 491770 453454
rect 492006 453218 522490 453454
rect 522726 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 399610 453134
rect 399846 452898 430330 453134
rect 430566 452898 461050 453134
rect 461286 452898 491770 453134
rect 492006 452898 522490 453134
rect 522726 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 40328 381454
rect 40564 381218 176056 381454
rect 176292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 220328 381454
rect 220564 381218 356056 381454
rect 356292 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 40328 381134
rect 40564 380898 176056 381134
rect 176292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 220328 381134
rect 220564 380898 356056 381134
rect 356292 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 41008 363454
rect 41244 363218 175376 363454
rect 175612 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 221008 363454
rect 221244 363218 355376 363454
rect 355612 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 41008 363134
rect 41244 362898 175376 363134
rect 175612 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 221008 363134
rect 221244 362898 355376 363134
rect 355612 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 40328 345454
rect 40564 345218 176056 345454
rect 176292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 40328 345134
rect 40564 344898 176056 345134
rect 176292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 41008 327454
rect 41244 327218 175376 327454
rect 175612 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 41008 327134
rect 41244 326898 175376 327134
rect 175612 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 40328 309454
rect 40564 309218 176056 309454
rect 176292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 40328 309134
rect 40564 308898 176056 309134
rect 176292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 114250 219454
rect 114486 219218 144970 219454
rect 145206 219218 175690 219454
rect 175926 219218 206410 219454
rect 206646 219218 237130 219454
rect 237366 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 114250 219134
rect 114486 218898 144970 219134
rect 145206 218898 175690 219134
rect 175926 218898 206410 219134
rect 206646 218898 237130 219134
rect 237366 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 129610 201454
rect 129846 201218 160330 201454
rect 160566 201218 191050 201454
rect 191286 201218 221770 201454
rect 222006 201218 252490 201454
rect 252726 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 129610 201134
rect 129846 200898 160330 201134
rect 160566 200898 191050 201134
rect 191286 200898 221770 201134
rect 222006 200898 252490 201134
rect 252726 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 114250 183454
rect 114486 183218 144970 183454
rect 145206 183218 175690 183454
rect 175926 183218 206410 183454
rect 206646 183218 237130 183454
rect 237366 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 114250 183134
rect 114486 182898 144970 183134
rect 145206 182898 175690 183134
rect 175926 182898 206410 183134
rect 206646 182898 237130 183134
rect 237366 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 129610 165454
rect 129846 165218 160330 165454
rect 160566 165218 191050 165454
rect 191286 165218 221770 165454
rect 222006 165218 252490 165454
rect 252726 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 129610 165134
rect 129846 164898 160330 165134
rect 160566 164898 191050 165134
rect 191286 164898 221770 165134
rect 222006 164898 252490 165134
rect 252726 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 264250 111454
rect 264486 111218 294970 111454
rect 295206 111218 325690 111454
rect 325926 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 264250 111134
rect 264486 110898 294970 111134
rect 295206 110898 325690 111134
rect 325926 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 279610 93454
rect 279846 93218 310330 93454
rect 310566 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 279610 93134
rect 279846 92898 310330 93134
rect 310566 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 264250 75454
rect 264486 75218 294970 75454
rect 295206 75218 325690 75454
rect 325926 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 264250 75134
rect 264486 74898 294970 75134
rect 295206 74898 325690 75134
rect 325926 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 279610 57454
rect 279846 57218 310330 57454
rect 310566 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 279610 57134
rect 279846 56898 310330 57134
rect 310566 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use merge_memory  merge_memory_inst
timestamp 0
transform 1 0 130000 0 1 460000
box 658 0 120000 39568
use sky130_sram_2kbyte_1rw1r_32x512_8  sky130_sram_2kbyte_1rw1r_32x512_8_inst0
timestamp 0
transform 1 0 220000 0 1 300000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sky130_sram_2kbyte_1rw1r_32x512_8_inst1
timestamp 0
transform 1 0 40000 0 1 300000
box 0 0 136620 83308
use wb_memory  wb_memory_inst
timestamp 0
transform 1 0 110000 0 1 160000
box 0 0 150000 70000
use wb_mux  wb_mux_inst
timestamp 0
transform 1 0 260000 0 1 40000
box 0 0 80000 79552
use wfg_top  wfg_top_inst
timestamp 0
transform 1 0 380000 0 1 440000
box 0 0 149210 110000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 158000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 158000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 158000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 158000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 158000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 232000 110414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 232000 146414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 232000 218414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 232000 254414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 122000 290414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 122000 326414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 385308 146414 458000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 232000 182414 458000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 385308 218414 458000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 385308 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 385308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 385308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 502000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 502000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 502000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 385308 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 385308 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 385308 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 552000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 552000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 552000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 552000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 158000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 158000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 158000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 158000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 122000 258134 158000 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 232000 114134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 232000 150134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 232000 222134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 232000 258134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 122000 294134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 122000 330134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 385308 150134 458000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 232000 186134 458000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 385308 222134 458000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 385308 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 385308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 385308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 502000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 502000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 502000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 385308 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 385308 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 385308 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 552000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 552000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 552000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 552000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 158000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 158000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 158000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 158000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 122000 261854 158000 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 232000 117854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 232000 153854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 232000 225854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 232000 261854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 122000 297854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 122000 333854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 385308 153854 458000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 232000 189854 458000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 385308 225854 458000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 385308 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 385308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 385308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 502000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 502000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 502000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 385308 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 385308 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 385308 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 552000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 552000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 552000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 552000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 158000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 158000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 158000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 158000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 232000 121574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 232000 157574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 232000 229574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 122000 265574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 122000 301574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 122000 337574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 385308 157574 458000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 232000 193574 458000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 385308 229574 458000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 385308 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 385308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 385308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 502000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 502000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 502000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 385308 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 385308 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 385308 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 552000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 552000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 552000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 552000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 232000 135854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 232000 171854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 232000 243854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 122000 279854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 122000 315854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 385308 135854 458000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 385308 171854 458000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 232000 207854 458000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 385308 243854 458000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 385308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 385308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 502000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 502000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 502000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 502000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 385308 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 385308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 385308 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 552000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 552000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 552000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 552000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 552000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 158000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 158000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 158000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 158000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 232000 139574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 232000 175574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 232000 247574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 122000 283574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 122000 319574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 438000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 438000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 438000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 438000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 385308 139574 458000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 385308 175574 458000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 232000 211574 458000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 385308 247574 458000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 385308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 385308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 502000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 502000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 502000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 502000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 385308 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 385308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 385308 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 552000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 552000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 552000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 552000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 232000 128414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 232000 164414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 232000 236414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 122000 272414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 122000 308414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 385308 128414 458000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 385308 164414 458000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 232000 200414 458000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 385308 236414 458000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 385308 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 385308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 502000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 502000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 502000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 502000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 385308 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 385308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 385308 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 552000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 552000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 552000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 552000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 552000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 232000 132134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 232000 168134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 232000 240134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 122000 276134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 122000 312134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 385308 132134 458000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 385308 168134 458000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 232000 204134 458000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 385308 240134 458000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 385308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 385308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 502000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 502000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 502000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 502000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 385308 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 385308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 385308 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 552000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 552000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 552000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 552000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 552000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
