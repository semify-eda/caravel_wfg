VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_mux
  CLASS BLOCK ;
  FOREIGN wb_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_ack_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.080 400.000 393.680 ;
    END
  END io_wbs_ack_0
  PIN io_wbs_ack_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END io_wbs_ack_1
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_adr_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1.400 400.000 2.000 ;
    END
  END io_wbs_adr_0[0]
  PIN io_wbs_adr_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.840 400.000 41.440 ;
    END
  END io_wbs_adr_0[10]
  PIN io_wbs_adr_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.920 400.000 45.520 ;
    END
  END io_wbs_adr_0[11]
  PIN io_wbs_adr_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 49.000 400.000 49.600 ;
    END
  END io_wbs_adr_0[12]
  PIN io_wbs_adr_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.080 400.000 53.680 ;
    END
  END io_wbs_adr_0[13]
  PIN io_wbs_adr_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.160 400.000 57.760 ;
    END
  END io_wbs_adr_0[14]
  PIN io_wbs_adr_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END io_wbs_adr_0[15]
  PIN io_wbs_adr_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 65.320 400.000 65.920 ;
    END
  END io_wbs_adr_0[16]
  PIN io_wbs_adr_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.720 400.000 69.320 ;
    END
  END io_wbs_adr_0[17]
  PIN io_wbs_adr_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.800 400.000 73.400 ;
    END
  END io_wbs_adr_0[18]
  PIN io_wbs_adr_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.880 400.000 77.480 ;
    END
  END io_wbs_adr_0[19]
  PIN io_wbs_adr_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.800 400.000 5.400 ;
    END
  END io_wbs_adr_0[1]
  PIN io_wbs_adr_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.960 400.000 81.560 ;
    END
  END io_wbs_adr_0[20]
  PIN io_wbs_adr_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END io_wbs_adr_0[21]
  PIN io_wbs_adr_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 89.120 400.000 89.720 ;
    END
  END io_wbs_adr_0[22]
  PIN io_wbs_adr_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 93.200 400.000 93.800 ;
    END
  END io_wbs_adr_0[23]
  PIN io_wbs_adr_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.280 400.000 97.880 ;
    END
  END io_wbs_adr_0[24]
  PIN io_wbs_adr_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 101.360 400.000 101.960 ;
    END
  END io_wbs_adr_0[25]
  PIN io_wbs_adr_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.760 400.000 105.360 ;
    END
  END io_wbs_adr_0[26]
  PIN io_wbs_adr_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END io_wbs_adr_0[27]
  PIN io_wbs_adr_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.920 400.000 113.520 ;
    END
  END io_wbs_adr_0[28]
  PIN io_wbs_adr_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.000 400.000 117.600 ;
    END
  END io_wbs_adr_0[29]
  PIN io_wbs_adr_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.880 400.000 9.480 ;
    END
  END io_wbs_adr_0[2]
  PIN io_wbs_adr_0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.080 400.000 121.680 ;
    END
  END io_wbs_adr_0[30]
  PIN io_wbs_adr_0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.160 400.000 125.760 ;
    END
  END io_wbs_adr_0[31]
  PIN io_wbs_adr_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 400.000 13.560 ;
    END
  END io_wbs_adr_0[3]
  PIN io_wbs_adr_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 400.000 17.640 ;
    END
  END io_wbs_adr_0[4]
  PIN io_wbs_adr_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.120 400.000 21.720 ;
    END
  END io_wbs_adr_0[5]
  PIN io_wbs_adr_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.200 400.000 25.800 ;
    END
  END io_wbs_adr_0[6]
  PIN io_wbs_adr_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.280 400.000 29.880 ;
    END
  END io_wbs_adr_0[7]
  PIN io_wbs_adr_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 33.360 400.000 33.960 ;
    END
  END io_wbs_adr_0[8]
  PIN io_wbs_adr_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.760 400.000 37.360 ;
    END
  END io_wbs_adr_0[9]
  PIN io_wbs_adr_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END io_wbs_adr_1[0]
  PIN io_wbs_adr_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_wbs_adr_1[10]
  PIN io_wbs_adr_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END io_wbs_adr_1[11]
  PIN io_wbs_adr_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_wbs_adr_1[12]
  PIN io_wbs_adr_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END io_wbs_adr_1[13]
  PIN io_wbs_adr_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_wbs_adr_1[14]
  PIN io_wbs_adr_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_wbs_adr_1[15]
  PIN io_wbs_adr_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END io_wbs_adr_1[16]
  PIN io_wbs_adr_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END io_wbs_adr_1[17]
  PIN io_wbs_adr_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END io_wbs_adr_1[18]
  PIN io_wbs_adr_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END io_wbs_adr_1[19]
  PIN io_wbs_adr_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_wbs_adr_1[1]
  PIN io_wbs_adr_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END io_wbs_adr_1[20]
  PIN io_wbs_adr_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_wbs_adr_1[21]
  PIN io_wbs_adr_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END io_wbs_adr_1[22]
  PIN io_wbs_adr_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END io_wbs_adr_1[23]
  PIN io_wbs_adr_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END io_wbs_adr_1[24]
  PIN io_wbs_adr_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END io_wbs_adr_1[25]
  PIN io_wbs_adr_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END io_wbs_adr_1[26]
  PIN io_wbs_adr_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_wbs_adr_1[27]
  PIN io_wbs_adr_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_wbs_adr_1[28]
  PIN io_wbs_adr_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_wbs_adr_1[29]
  PIN io_wbs_adr_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_wbs_adr_1[2]
  PIN io_wbs_adr_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END io_wbs_adr_1[30]
  PIN io_wbs_adr_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END io_wbs_adr_1[31]
  PIN io_wbs_adr_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END io_wbs_adr_1[3]
  PIN io_wbs_adr_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_wbs_adr_1[4]
  PIN io_wbs_adr_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_wbs_adr_1[5]
  PIN io_wbs_adr_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END io_wbs_adr_1[6]
  PIN io_wbs_adr_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END io_wbs_adr_1[7]
  PIN io_wbs_adr_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_wbs_adr_1[8]
  PIN io_wbs_adr_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END io_wbs_adr_1[9]
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_cyc_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END io_wbs_cyc_0
  PIN io_wbs_cyc_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END io_wbs_cyc_1
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datrd_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.080 400.000 257.680 ;
    END
  END io_wbs_datrd_0[0]
  PIN io_wbs_datrd_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.200 400.000 297.800 ;
    END
  END io_wbs_datrd_0[10]
  PIN io_wbs_datrd_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.280 400.000 301.880 ;
    END
  END io_wbs_datrd_0[11]
  PIN io_wbs_datrd_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.680 400.000 305.280 ;
    END
  END io_wbs_datrd_0[12]
  PIN io_wbs_datrd_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.760 400.000 309.360 ;
    END
  END io_wbs_datrd_0[13]
  PIN io_wbs_datrd_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.840 400.000 313.440 ;
    END
  END io_wbs_datrd_0[14]
  PIN io_wbs_datrd_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.920 400.000 317.520 ;
    END
  END io_wbs_datrd_0[15]
  PIN io_wbs_datrd_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END io_wbs_datrd_0[16]
  PIN io_wbs_datrd_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.080 400.000 325.680 ;
    END
  END io_wbs_datrd_0[17]
  PIN io_wbs_datrd_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.160 400.000 329.760 ;
    END
  END io_wbs_datrd_0[18]
  PIN io_wbs_datrd_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.240 400.000 333.840 ;
    END
  END io_wbs_datrd_0[19]
  PIN io_wbs_datrd_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.160 400.000 261.760 ;
    END
  END io_wbs_datrd_0[1]
  PIN io_wbs_datrd_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 336.640 400.000 337.240 ;
    END
  END io_wbs_datrd_0[20]
  PIN io_wbs_datrd_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.720 400.000 341.320 ;
    END
  END io_wbs_datrd_0[21]
  PIN io_wbs_datrd_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.800 400.000 345.400 ;
    END
  END io_wbs_datrd_0[22]
  PIN io_wbs_datrd_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.880 400.000 349.480 ;
    END
  END io_wbs_datrd_0[23]
  PIN io_wbs_datrd_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.960 400.000 353.560 ;
    END
  END io_wbs_datrd_0[24]
  PIN io_wbs_datrd_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.040 400.000 357.640 ;
    END
  END io_wbs_datrd_0[25]
  PIN io_wbs_datrd_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END io_wbs_datrd_0[26]
  PIN io_wbs_datrd_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.200 400.000 365.800 ;
    END
  END io_wbs_datrd_0[27]
  PIN io_wbs_datrd_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 368.600 400.000 369.200 ;
    END
  END io_wbs_datrd_0[28]
  PIN io_wbs_datrd_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END io_wbs_datrd_0[29]
  PIN io_wbs_datrd_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END io_wbs_datrd_0[2]
  PIN io_wbs_datrd_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.760 400.000 377.360 ;
    END
  END io_wbs_datrd_0[30]
  PIN io_wbs_datrd_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END io_wbs_datrd_0[31]
  PIN io_wbs_datrd_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END io_wbs_datrd_0[3]
  PIN io_wbs_datrd_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.720 400.000 273.320 ;
    END
  END io_wbs_datrd_0[4]
  PIN io_wbs_datrd_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.800 400.000 277.400 ;
    END
  END io_wbs_datrd_0[5]
  PIN io_wbs_datrd_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.880 400.000 281.480 ;
    END
  END io_wbs_datrd_0[6]
  PIN io_wbs_datrd_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.960 400.000 285.560 ;
    END
  END io_wbs_datrd_0[7]
  PIN io_wbs_datrd_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.040 400.000 289.640 ;
    END
  END io_wbs_datrd_0[8]
  PIN io_wbs_datrd_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END io_wbs_datrd_0[9]
  PIN io_wbs_datrd_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_wbs_datrd_1[0]
  PIN io_wbs_datrd_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END io_wbs_datrd_1[10]
  PIN io_wbs_datrd_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END io_wbs_datrd_1[11]
  PIN io_wbs_datrd_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END io_wbs_datrd_1[12]
  PIN io_wbs_datrd_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END io_wbs_datrd_1[13]
  PIN io_wbs_datrd_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END io_wbs_datrd_1[14]
  PIN io_wbs_datrd_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END io_wbs_datrd_1[15]
  PIN io_wbs_datrd_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END io_wbs_datrd_1[16]
  PIN io_wbs_datrd_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END io_wbs_datrd_1[17]
  PIN io_wbs_datrd_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END io_wbs_datrd_1[18]
  PIN io_wbs_datrd_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_wbs_datrd_1[19]
  PIN io_wbs_datrd_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END io_wbs_datrd_1[1]
  PIN io_wbs_datrd_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END io_wbs_datrd_1[20]
  PIN io_wbs_datrd_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END io_wbs_datrd_1[21]
  PIN io_wbs_datrd_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END io_wbs_datrd_1[22]
  PIN io_wbs_datrd_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END io_wbs_datrd_1[23]
  PIN io_wbs_datrd_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END io_wbs_datrd_1[24]
  PIN io_wbs_datrd_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END io_wbs_datrd_1[25]
  PIN io_wbs_datrd_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END io_wbs_datrd_1[26]
  PIN io_wbs_datrd_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END io_wbs_datrd_1[27]
  PIN io_wbs_datrd_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END io_wbs_datrd_1[28]
  PIN io_wbs_datrd_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END io_wbs_datrd_1[29]
  PIN io_wbs_datrd_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_wbs_datrd_1[2]
  PIN io_wbs_datrd_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_wbs_datrd_1[30]
  PIN io_wbs_datrd_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_wbs_datrd_1[31]
  PIN io_wbs_datrd_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END io_wbs_datrd_1[3]
  PIN io_wbs_datrd_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END io_wbs_datrd_1[4]
  PIN io_wbs_datrd_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END io_wbs_datrd_1[5]
  PIN io_wbs_datrd_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END io_wbs_datrd_1[6]
  PIN io_wbs_datrd_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END io_wbs_datrd_1[7]
  PIN io_wbs_datrd_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_wbs_datrd_1[8]
  PIN io_wbs_datrd_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END io_wbs_datrd_1[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_datwr_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END io_wbs_datwr_0[0]
  PIN io_wbs_datwr_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.680 400.000 169.280 ;
    END
  END io_wbs_datwr_0[10]
  PIN io_wbs_datwr_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.760 400.000 173.360 ;
    END
  END io_wbs_datwr_0[11]
  PIN io_wbs_datwr_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END io_wbs_datwr_0[12]
  PIN io_wbs_datwr_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.920 400.000 181.520 ;
    END
  END io_wbs_datwr_0[13]
  PIN io_wbs_datwr_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 185.000 400.000 185.600 ;
    END
  END io_wbs_datwr_0[14]
  PIN io_wbs_datwr_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END io_wbs_datwr_0[15]
  PIN io_wbs_datwr_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.160 400.000 193.760 ;
    END
  END io_wbs_datwr_0[16]
  PIN io_wbs_datwr_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END io_wbs_datwr_0[17]
  PIN io_wbs_datwr_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 201.320 400.000 201.920 ;
    END
  END io_wbs_datwr_0[18]
  PIN io_wbs_datwr_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 400.000 205.320 ;
    END
  END io_wbs_datwr_0[19]
  PIN io_wbs_datwr_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 133.320 400.000 133.920 ;
    END
  END io_wbs_datwr_0[1]
  PIN io_wbs_datwr_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.800 400.000 209.400 ;
    END
  END io_wbs_datwr_0[20]
  PIN io_wbs_datwr_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 400.000 213.480 ;
    END
  END io_wbs_datwr_0[21]
  PIN io_wbs_datwr_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 400.000 217.560 ;
    END
  END io_wbs_datwr_0[22]
  PIN io_wbs_datwr_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 400.000 221.640 ;
    END
  END io_wbs_datwr_0[23]
  PIN io_wbs_datwr_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.120 400.000 225.720 ;
    END
  END io_wbs_datwr_0[24]
  PIN io_wbs_datwr_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.200 400.000 229.800 ;
    END
  END io_wbs_datwr_0[25]
  PIN io_wbs_datwr_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.280 400.000 233.880 ;
    END
  END io_wbs_datwr_0[26]
  PIN io_wbs_datwr_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.680 400.000 237.280 ;
    END
  END io_wbs_datwr_0[27]
  PIN io_wbs_datwr_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.760 400.000 241.360 ;
    END
  END io_wbs_datwr_0[28]
  PIN io_wbs_datwr_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.840 400.000 245.440 ;
    END
  END io_wbs_datwr_0[29]
  PIN io_wbs_datwr_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.720 400.000 137.320 ;
    END
  END io_wbs_datwr_0[2]
  PIN io_wbs_datwr_0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.920 400.000 249.520 ;
    END
  END io_wbs_datwr_0[30]
  PIN io_wbs_datwr_0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.000 400.000 253.600 ;
    END
  END io_wbs_datwr_0[31]
  PIN io_wbs_datwr_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.800 400.000 141.400 ;
    END
  END io_wbs_datwr_0[3]
  PIN io_wbs_datwr_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.880 400.000 145.480 ;
    END
  END io_wbs_datwr_0[4]
  PIN io_wbs_datwr_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.960 400.000 149.560 ;
    END
  END io_wbs_datwr_0[5]
  PIN io_wbs_datwr_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 400.000 153.640 ;
    END
  END io_wbs_datwr_0[6]
  PIN io_wbs_datwr_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.120 400.000 157.720 ;
    END
  END io_wbs_datwr_0[7]
  PIN io_wbs_datwr_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.200 400.000 161.800 ;
    END
  END io_wbs_datwr_0[8]
  PIN io_wbs_datwr_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.280 400.000 165.880 ;
    END
  END io_wbs_datwr_0[9]
  PIN io_wbs_datwr_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_wbs_datwr_1[0]
  PIN io_wbs_datwr_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END io_wbs_datwr_1[10]
  PIN io_wbs_datwr_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_wbs_datwr_1[11]
  PIN io_wbs_datwr_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_wbs_datwr_1[12]
  PIN io_wbs_datwr_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END io_wbs_datwr_1[13]
  PIN io_wbs_datwr_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END io_wbs_datwr_1[14]
  PIN io_wbs_datwr_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END io_wbs_datwr_1[15]
  PIN io_wbs_datwr_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_wbs_datwr_1[16]
  PIN io_wbs_datwr_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_wbs_datwr_1[17]
  PIN io_wbs_datwr_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END io_wbs_datwr_1[18]
  PIN io_wbs_datwr_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_wbs_datwr_1[19]
  PIN io_wbs_datwr_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_wbs_datwr_1[1]
  PIN io_wbs_datwr_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END io_wbs_datwr_1[20]
  PIN io_wbs_datwr_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END io_wbs_datwr_1[21]
  PIN io_wbs_datwr_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_wbs_datwr_1[22]
  PIN io_wbs_datwr_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_wbs_datwr_1[23]
  PIN io_wbs_datwr_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END io_wbs_datwr_1[24]
  PIN io_wbs_datwr_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_wbs_datwr_1[25]
  PIN io_wbs_datwr_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END io_wbs_datwr_1[26]
  PIN io_wbs_datwr_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_wbs_datwr_1[27]
  PIN io_wbs_datwr_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END io_wbs_datwr_1[28]
  PIN io_wbs_datwr_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_wbs_datwr_1[29]
  PIN io_wbs_datwr_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END io_wbs_datwr_1[2]
  PIN io_wbs_datwr_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_wbs_datwr_1[30]
  PIN io_wbs_datwr_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_wbs_datwr_1[31]
  PIN io_wbs_datwr_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END io_wbs_datwr_1[3]
  PIN io_wbs_datwr_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END io_wbs_datwr_1[4]
  PIN io_wbs_datwr_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END io_wbs_datwr_1[5]
  PIN io_wbs_datwr_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_wbs_datwr_1[6]
  PIN io_wbs_datwr_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END io_wbs_datwr_1[7]
  PIN io_wbs_datwr_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END io_wbs_datwr_1[8]
  PIN io_wbs_datwr_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END io_wbs_datwr_1[9]
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_stb_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END io_wbs_stb_0
  PIN io_wbs_stb_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END io_wbs_stb_1
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END io_wbs_we
  PIN io_wbs_we_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.920 400.000 385.520 ;
    END
  END io_wbs_we_0
  PIN io_wbs_we_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END io_wbs_we_1
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 1.910 8.540 398.290 389.200 ;
      LAYER met2 ;
        RECT 1.940 4.280 398.260 397.645 ;
        RECT 2.490 1.515 5.330 4.280 ;
        RECT 6.170 1.515 9.470 4.280 ;
        RECT 10.310 1.515 13.610 4.280 ;
        RECT 14.450 1.515 17.290 4.280 ;
        RECT 18.130 1.515 21.430 4.280 ;
        RECT 22.270 1.515 25.570 4.280 ;
        RECT 26.410 1.515 29.250 4.280 ;
        RECT 30.090 1.515 33.390 4.280 ;
        RECT 34.230 1.515 37.530 4.280 ;
        RECT 38.370 1.515 41.670 4.280 ;
        RECT 42.510 1.515 45.350 4.280 ;
        RECT 46.190 1.515 49.490 4.280 ;
        RECT 50.330 1.515 53.630 4.280 ;
        RECT 54.470 1.515 57.310 4.280 ;
        RECT 58.150 1.515 61.450 4.280 ;
        RECT 62.290 1.515 65.590 4.280 ;
        RECT 66.430 1.515 69.270 4.280 ;
        RECT 70.110 1.515 73.410 4.280 ;
        RECT 74.250 1.515 77.550 4.280 ;
        RECT 78.390 1.515 81.690 4.280 ;
        RECT 82.530 1.515 85.370 4.280 ;
        RECT 86.210 1.515 89.510 4.280 ;
        RECT 90.350 1.515 93.650 4.280 ;
        RECT 94.490 1.515 97.330 4.280 ;
        RECT 98.170 1.515 101.470 4.280 ;
        RECT 102.310 1.515 105.610 4.280 ;
        RECT 106.450 1.515 109.290 4.280 ;
        RECT 110.130 1.515 113.430 4.280 ;
        RECT 114.270 1.515 117.570 4.280 ;
        RECT 118.410 1.515 121.710 4.280 ;
        RECT 122.550 1.515 125.390 4.280 ;
        RECT 126.230 1.515 129.530 4.280 ;
        RECT 130.370 1.515 133.670 4.280 ;
        RECT 134.510 1.515 137.350 4.280 ;
        RECT 138.190 1.515 141.490 4.280 ;
        RECT 142.330 1.515 145.630 4.280 ;
        RECT 146.470 1.515 149.310 4.280 ;
        RECT 150.150 1.515 153.450 4.280 ;
        RECT 154.290 1.515 157.590 4.280 ;
        RECT 158.430 1.515 161.730 4.280 ;
        RECT 162.570 1.515 165.410 4.280 ;
        RECT 166.250 1.515 169.550 4.280 ;
        RECT 170.390 1.515 173.690 4.280 ;
        RECT 174.530 1.515 177.370 4.280 ;
        RECT 178.210 1.515 181.510 4.280 ;
        RECT 182.350 1.515 185.650 4.280 ;
        RECT 186.490 1.515 189.330 4.280 ;
        RECT 190.170 1.515 193.470 4.280 ;
        RECT 194.310 1.515 197.610 4.280 ;
        RECT 198.450 1.515 201.750 4.280 ;
        RECT 202.590 1.515 205.430 4.280 ;
        RECT 206.270 1.515 209.570 4.280 ;
        RECT 210.410 1.515 213.710 4.280 ;
        RECT 214.550 1.515 217.390 4.280 ;
        RECT 218.230 1.515 221.530 4.280 ;
        RECT 222.370 1.515 225.670 4.280 ;
        RECT 226.510 1.515 229.350 4.280 ;
        RECT 230.190 1.515 233.490 4.280 ;
        RECT 234.330 1.515 237.630 4.280 ;
        RECT 238.470 1.515 241.770 4.280 ;
        RECT 242.610 1.515 245.450 4.280 ;
        RECT 246.290 1.515 249.590 4.280 ;
        RECT 250.430 1.515 253.730 4.280 ;
        RECT 254.570 1.515 257.410 4.280 ;
        RECT 258.250 1.515 261.550 4.280 ;
        RECT 262.390 1.515 265.690 4.280 ;
        RECT 266.530 1.515 269.370 4.280 ;
        RECT 270.210 1.515 273.510 4.280 ;
        RECT 274.350 1.515 277.650 4.280 ;
        RECT 278.490 1.515 281.790 4.280 ;
        RECT 282.630 1.515 285.470 4.280 ;
        RECT 286.310 1.515 289.610 4.280 ;
        RECT 290.450 1.515 293.750 4.280 ;
        RECT 294.590 1.515 297.430 4.280 ;
        RECT 298.270 1.515 301.570 4.280 ;
        RECT 302.410 1.515 305.710 4.280 ;
        RECT 306.550 1.515 309.390 4.280 ;
        RECT 310.230 1.515 313.530 4.280 ;
        RECT 314.370 1.515 317.670 4.280 ;
        RECT 318.510 1.515 321.810 4.280 ;
        RECT 322.650 1.515 325.490 4.280 ;
        RECT 326.330 1.515 329.630 4.280 ;
        RECT 330.470 1.515 333.770 4.280 ;
        RECT 334.610 1.515 337.450 4.280 ;
        RECT 338.290 1.515 341.590 4.280 ;
        RECT 342.430 1.515 345.730 4.280 ;
        RECT 346.570 1.515 349.410 4.280 ;
        RECT 350.250 1.515 353.550 4.280 ;
        RECT 354.390 1.515 357.690 4.280 ;
        RECT 358.530 1.515 361.830 4.280 ;
        RECT 362.670 1.515 365.510 4.280 ;
        RECT 366.350 1.515 369.650 4.280 ;
        RECT 370.490 1.515 373.790 4.280 ;
        RECT 374.630 1.515 377.470 4.280 ;
        RECT 378.310 1.515 381.610 4.280 ;
        RECT 382.450 1.515 385.750 4.280 ;
        RECT 386.590 1.515 389.430 4.280 ;
        RECT 390.270 1.515 393.570 4.280 ;
        RECT 394.410 1.515 397.710 4.280 ;
      LAYER met3 ;
        RECT 4.400 396.760 395.600 397.625 ;
        RECT 4.000 394.080 396.000 396.760 ;
        RECT 4.400 392.680 395.600 394.080 ;
        RECT 4.000 390.000 396.000 392.680 ;
        RECT 4.400 388.600 395.600 390.000 ;
        RECT 4.000 385.920 396.000 388.600 ;
        RECT 4.400 384.520 395.600 385.920 ;
        RECT 4.000 381.840 396.000 384.520 ;
        RECT 4.400 380.440 395.600 381.840 ;
        RECT 4.000 377.760 396.000 380.440 ;
        RECT 4.400 376.360 395.600 377.760 ;
        RECT 4.000 373.680 396.000 376.360 ;
        RECT 4.400 372.280 395.600 373.680 ;
        RECT 4.000 369.600 396.000 372.280 ;
        RECT 4.400 368.200 395.600 369.600 ;
        RECT 4.000 366.200 396.000 368.200 ;
        RECT 4.400 364.800 395.600 366.200 ;
        RECT 4.000 362.120 396.000 364.800 ;
        RECT 4.400 360.720 395.600 362.120 ;
        RECT 4.000 358.040 396.000 360.720 ;
        RECT 4.400 356.640 395.600 358.040 ;
        RECT 4.000 353.960 396.000 356.640 ;
        RECT 4.400 352.560 395.600 353.960 ;
        RECT 4.000 349.880 396.000 352.560 ;
        RECT 4.400 348.480 395.600 349.880 ;
        RECT 4.000 345.800 396.000 348.480 ;
        RECT 4.400 344.400 395.600 345.800 ;
        RECT 4.000 341.720 396.000 344.400 ;
        RECT 4.400 340.320 395.600 341.720 ;
        RECT 4.000 337.640 396.000 340.320 ;
        RECT 4.400 336.240 395.600 337.640 ;
        RECT 4.000 334.240 396.000 336.240 ;
        RECT 4.400 332.840 395.600 334.240 ;
        RECT 4.000 330.160 396.000 332.840 ;
        RECT 4.400 328.760 395.600 330.160 ;
        RECT 4.000 326.080 396.000 328.760 ;
        RECT 4.400 324.680 395.600 326.080 ;
        RECT 4.000 322.000 396.000 324.680 ;
        RECT 4.400 320.600 395.600 322.000 ;
        RECT 4.000 317.920 396.000 320.600 ;
        RECT 4.400 316.520 395.600 317.920 ;
        RECT 4.000 313.840 396.000 316.520 ;
        RECT 4.400 312.440 395.600 313.840 ;
        RECT 4.000 309.760 396.000 312.440 ;
        RECT 4.400 308.360 395.600 309.760 ;
        RECT 4.000 305.680 396.000 308.360 ;
        RECT 4.400 304.280 395.600 305.680 ;
        RECT 4.000 302.280 396.000 304.280 ;
        RECT 4.400 300.880 395.600 302.280 ;
        RECT 4.000 298.200 396.000 300.880 ;
        RECT 4.400 296.800 395.600 298.200 ;
        RECT 4.000 294.120 396.000 296.800 ;
        RECT 4.400 292.720 395.600 294.120 ;
        RECT 4.000 290.040 396.000 292.720 ;
        RECT 4.400 288.640 395.600 290.040 ;
        RECT 4.000 285.960 396.000 288.640 ;
        RECT 4.400 284.560 395.600 285.960 ;
        RECT 4.000 281.880 396.000 284.560 ;
        RECT 4.400 280.480 395.600 281.880 ;
        RECT 4.000 277.800 396.000 280.480 ;
        RECT 4.400 276.400 395.600 277.800 ;
        RECT 4.000 273.720 396.000 276.400 ;
        RECT 4.400 272.320 395.600 273.720 ;
        RECT 4.000 269.640 396.000 272.320 ;
        RECT 4.400 268.240 395.600 269.640 ;
        RECT 4.000 266.240 396.000 268.240 ;
        RECT 4.400 264.840 395.600 266.240 ;
        RECT 4.000 262.160 396.000 264.840 ;
        RECT 4.400 260.760 395.600 262.160 ;
        RECT 4.000 258.080 396.000 260.760 ;
        RECT 4.400 256.680 395.600 258.080 ;
        RECT 4.000 254.000 396.000 256.680 ;
        RECT 4.400 252.600 395.600 254.000 ;
        RECT 4.000 249.920 396.000 252.600 ;
        RECT 4.400 248.520 395.600 249.920 ;
        RECT 4.000 245.840 396.000 248.520 ;
        RECT 4.400 244.440 395.600 245.840 ;
        RECT 4.000 241.760 396.000 244.440 ;
        RECT 4.400 240.360 395.600 241.760 ;
        RECT 4.000 237.680 396.000 240.360 ;
        RECT 4.400 236.280 395.600 237.680 ;
        RECT 4.000 234.280 396.000 236.280 ;
        RECT 4.400 232.880 395.600 234.280 ;
        RECT 4.000 230.200 396.000 232.880 ;
        RECT 4.400 228.800 395.600 230.200 ;
        RECT 4.000 226.120 396.000 228.800 ;
        RECT 4.400 224.720 395.600 226.120 ;
        RECT 4.000 222.040 396.000 224.720 ;
        RECT 4.400 220.640 395.600 222.040 ;
        RECT 4.000 217.960 396.000 220.640 ;
        RECT 4.400 216.560 395.600 217.960 ;
        RECT 4.000 213.880 396.000 216.560 ;
        RECT 4.400 212.480 395.600 213.880 ;
        RECT 4.000 209.800 396.000 212.480 ;
        RECT 4.400 208.400 395.600 209.800 ;
        RECT 4.000 205.720 396.000 208.400 ;
        RECT 4.400 204.320 395.600 205.720 ;
        RECT 4.000 202.320 396.000 204.320 ;
        RECT 4.400 200.920 395.600 202.320 ;
        RECT 4.000 198.240 396.000 200.920 ;
        RECT 4.400 196.840 395.600 198.240 ;
        RECT 4.000 194.160 396.000 196.840 ;
        RECT 4.400 192.760 395.600 194.160 ;
        RECT 4.000 190.080 396.000 192.760 ;
        RECT 4.400 188.680 395.600 190.080 ;
        RECT 4.000 186.000 396.000 188.680 ;
        RECT 4.400 184.600 395.600 186.000 ;
        RECT 4.000 181.920 396.000 184.600 ;
        RECT 4.400 180.520 395.600 181.920 ;
        RECT 4.000 177.840 396.000 180.520 ;
        RECT 4.400 176.440 395.600 177.840 ;
        RECT 4.000 173.760 396.000 176.440 ;
        RECT 4.400 172.360 395.600 173.760 ;
        RECT 4.000 169.680 396.000 172.360 ;
        RECT 4.400 168.280 395.600 169.680 ;
        RECT 4.000 166.280 396.000 168.280 ;
        RECT 4.400 164.880 395.600 166.280 ;
        RECT 4.000 162.200 396.000 164.880 ;
        RECT 4.400 160.800 395.600 162.200 ;
        RECT 4.000 158.120 396.000 160.800 ;
        RECT 4.400 156.720 395.600 158.120 ;
        RECT 4.000 154.040 396.000 156.720 ;
        RECT 4.400 152.640 395.600 154.040 ;
        RECT 4.000 149.960 396.000 152.640 ;
        RECT 4.400 148.560 395.600 149.960 ;
        RECT 4.000 145.880 396.000 148.560 ;
        RECT 4.400 144.480 395.600 145.880 ;
        RECT 4.000 141.800 396.000 144.480 ;
        RECT 4.400 140.400 395.600 141.800 ;
        RECT 4.000 137.720 396.000 140.400 ;
        RECT 4.400 136.320 395.600 137.720 ;
        RECT 4.000 134.320 396.000 136.320 ;
        RECT 4.400 132.920 395.600 134.320 ;
        RECT 4.000 130.240 396.000 132.920 ;
        RECT 4.400 128.840 395.600 130.240 ;
        RECT 4.000 126.160 396.000 128.840 ;
        RECT 4.400 124.760 395.600 126.160 ;
        RECT 4.000 122.080 396.000 124.760 ;
        RECT 4.400 120.680 395.600 122.080 ;
        RECT 4.000 118.000 396.000 120.680 ;
        RECT 4.400 116.600 395.600 118.000 ;
        RECT 4.000 113.920 396.000 116.600 ;
        RECT 4.400 112.520 395.600 113.920 ;
        RECT 4.000 109.840 396.000 112.520 ;
        RECT 4.400 108.440 395.600 109.840 ;
        RECT 4.000 105.760 396.000 108.440 ;
        RECT 4.400 104.360 395.600 105.760 ;
        RECT 4.000 102.360 396.000 104.360 ;
        RECT 4.400 100.960 395.600 102.360 ;
        RECT 4.000 98.280 396.000 100.960 ;
        RECT 4.400 96.880 395.600 98.280 ;
        RECT 4.000 94.200 396.000 96.880 ;
        RECT 4.400 92.800 395.600 94.200 ;
        RECT 4.000 90.120 396.000 92.800 ;
        RECT 4.400 88.720 395.600 90.120 ;
        RECT 4.000 86.040 396.000 88.720 ;
        RECT 4.400 84.640 395.600 86.040 ;
        RECT 4.000 81.960 396.000 84.640 ;
        RECT 4.400 80.560 395.600 81.960 ;
        RECT 4.000 77.880 396.000 80.560 ;
        RECT 4.400 76.480 395.600 77.880 ;
        RECT 4.000 73.800 396.000 76.480 ;
        RECT 4.400 72.400 395.600 73.800 ;
        RECT 4.000 69.720 396.000 72.400 ;
        RECT 4.400 68.320 395.600 69.720 ;
        RECT 4.000 66.320 396.000 68.320 ;
        RECT 4.400 64.920 395.600 66.320 ;
        RECT 4.000 62.240 396.000 64.920 ;
        RECT 4.400 60.840 395.600 62.240 ;
        RECT 4.000 58.160 396.000 60.840 ;
        RECT 4.400 56.760 395.600 58.160 ;
        RECT 4.000 54.080 396.000 56.760 ;
        RECT 4.400 52.680 395.600 54.080 ;
        RECT 4.000 50.000 396.000 52.680 ;
        RECT 4.400 48.600 395.600 50.000 ;
        RECT 4.000 45.920 396.000 48.600 ;
        RECT 4.400 44.520 395.600 45.920 ;
        RECT 4.000 41.840 396.000 44.520 ;
        RECT 4.400 40.440 395.600 41.840 ;
        RECT 4.000 37.760 396.000 40.440 ;
        RECT 4.400 36.360 395.600 37.760 ;
        RECT 4.000 34.360 396.000 36.360 ;
        RECT 4.400 32.960 395.600 34.360 ;
        RECT 4.000 30.280 396.000 32.960 ;
        RECT 4.400 28.880 395.600 30.280 ;
        RECT 4.000 26.200 396.000 28.880 ;
        RECT 4.400 24.800 395.600 26.200 ;
        RECT 4.000 22.120 396.000 24.800 ;
        RECT 4.400 20.720 395.600 22.120 ;
        RECT 4.000 18.040 396.000 20.720 ;
        RECT 4.400 16.640 395.600 18.040 ;
        RECT 4.000 13.960 396.000 16.640 ;
        RECT 4.400 12.560 395.600 13.960 ;
        RECT 4.000 9.880 396.000 12.560 ;
        RECT 4.400 8.480 395.600 9.880 ;
        RECT 4.000 5.800 396.000 8.480 ;
        RECT 4.400 4.400 395.600 5.800 ;
        RECT 4.000 2.400 396.000 4.400 ;
        RECT 4.400 1.535 395.600 2.400 ;
  END
END wb_mux
END LIBRARY

