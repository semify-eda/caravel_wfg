magic
tech sky130A
magscale 1 2
timestamp 1656942120
<< obsli1 >>
rect 1104 2159 118864 67473
<< obsm1 >>
rect 566 8 119402 67584
<< metal2 >>
rect 1306 69200 1362 70000
rect 3882 69200 3938 70000
rect 6458 69200 6514 70000
rect 9126 69200 9182 70000
rect 11702 69200 11758 70000
rect 14278 69200 14334 70000
rect 16946 69200 17002 70000
rect 19522 69200 19578 70000
rect 22098 69200 22154 70000
rect 24766 69200 24822 70000
rect 27342 69200 27398 70000
rect 29918 69200 29974 70000
rect 32586 69200 32642 70000
rect 35162 69200 35218 70000
rect 37738 69200 37794 70000
rect 40406 69200 40462 70000
rect 42982 69200 43038 70000
rect 45558 69200 45614 70000
rect 48226 69200 48282 70000
rect 50802 69200 50858 70000
rect 53378 69200 53434 70000
rect 56046 69200 56102 70000
rect 58622 69200 58678 70000
rect 61290 69200 61346 70000
rect 63866 69200 63922 70000
rect 66442 69200 66498 70000
rect 69110 69200 69166 70000
rect 71686 69200 71742 70000
rect 74262 69200 74318 70000
rect 76930 69200 76986 70000
rect 79506 69200 79562 70000
rect 82082 69200 82138 70000
rect 84750 69200 84806 70000
rect 87326 69200 87382 70000
rect 89902 69200 89958 70000
rect 92570 69200 92626 70000
rect 95146 69200 95202 70000
rect 97722 69200 97778 70000
rect 100390 69200 100446 70000
rect 102966 69200 103022 70000
rect 105542 69200 105598 70000
rect 108210 69200 108266 70000
rect 110786 69200 110842 70000
rect 113362 69200 113418 70000
rect 116030 69200 116086 70000
rect 118606 69200 118662 70000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5262 0 5318 800
rect 6366 0 6422 800
rect 7562 0 7618 800
rect 8758 0 8814 800
rect 9954 0 10010 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13450 0 13506 800
rect 14646 0 14702 800
rect 15842 0 15898 800
rect 16946 0 17002 800
rect 18142 0 18198 800
rect 19338 0 19394 800
rect 20534 0 20590 800
rect 21730 0 21786 800
rect 22834 0 22890 800
rect 24030 0 24086 800
rect 25226 0 25282 800
rect 26422 0 26478 800
rect 27618 0 27674 800
rect 28722 0 28778 800
rect 29918 0 29974 800
rect 31114 0 31170 800
rect 32310 0 32366 800
rect 33414 0 33470 800
rect 34610 0 34666 800
rect 35806 0 35862 800
rect 37002 0 37058 800
rect 38198 0 38254 800
rect 39302 0 39358 800
rect 40498 0 40554 800
rect 41694 0 41750 800
rect 42890 0 42946 800
rect 44086 0 44142 800
rect 45190 0 45246 800
rect 46386 0 46442 800
rect 47582 0 47638 800
rect 48778 0 48834 800
rect 49882 0 49938 800
rect 51078 0 51134 800
rect 52274 0 52330 800
rect 53470 0 53526 800
rect 54666 0 54722 800
rect 55770 0 55826 800
rect 56966 0 57022 800
rect 58162 0 58218 800
rect 59358 0 59414 800
rect 60554 0 60610 800
rect 61658 0 61714 800
rect 62854 0 62910 800
rect 64050 0 64106 800
rect 65246 0 65302 800
rect 66350 0 66406 800
rect 67546 0 67602 800
rect 68742 0 68798 800
rect 69938 0 69994 800
rect 71134 0 71190 800
rect 72238 0 72294 800
rect 73434 0 73490 800
rect 74630 0 74686 800
rect 75826 0 75882 800
rect 76930 0 76986 800
rect 78126 0 78182 800
rect 79322 0 79378 800
rect 80518 0 80574 800
rect 81714 0 81770 800
rect 82818 0 82874 800
rect 84014 0 84070 800
rect 85210 0 85266 800
rect 86406 0 86462 800
rect 87602 0 87658 800
rect 88706 0 88762 800
rect 89902 0 89958 800
rect 91098 0 91154 800
rect 92294 0 92350 800
rect 93398 0 93454 800
rect 94594 0 94650 800
rect 95790 0 95846 800
rect 96986 0 97042 800
rect 98182 0 98238 800
rect 99286 0 99342 800
rect 100482 0 100538 800
rect 101678 0 101734 800
rect 102874 0 102930 800
rect 104070 0 104126 800
rect 105174 0 105230 800
rect 106370 0 106426 800
rect 107566 0 107622 800
rect 108762 0 108818 800
rect 109866 0 109922 800
rect 111062 0 111118 800
rect 112258 0 112314 800
rect 113454 0 113510 800
rect 114650 0 114706 800
rect 115754 0 115810 800
rect 116950 0 117006 800
rect 118146 0 118202 800
rect 119342 0 119398 800
<< obsm2 >>
rect 572 69144 1250 69306
rect 1418 69144 3826 69306
rect 3994 69144 6402 69306
rect 6570 69144 9070 69306
rect 9238 69144 11646 69306
rect 11814 69144 14222 69306
rect 14390 69144 16890 69306
rect 17058 69144 19466 69306
rect 19634 69144 22042 69306
rect 22210 69144 24710 69306
rect 24878 69144 27286 69306
rect 27454 69144 29862 69306
rect 30030 69144 32530 69306
rect 32698 69144 35106 69306
rect 35274 69144 37682 69306
rect 37850 69144 40350 69306
rect 40518 69144 42926 69306
rect 43094 69144 45502 69306
rect 45670 69144 48170 69306
rect 48338 69144 50746 69306
rect 50914 69144 53322 69306
rect 53490 69144 55990 69306
rect 56158 69144 58566 69306
rect 58734 69144 61234 69306
rect 61402 69144 63810 69306
rect 63978 69144 66386 69306
rect 66554 69144 69054 69306
rect 69222 69144 71630 69306
rect 71798 69144 74206 69306
rect 74374 69144 76874 69306
rect 77042 69144 79450 69306
rect 79618 69144 82026 69306
rect 82194 69144 84694 69306
rect 84862 69144 87270 69306
rect 87438 69144 89846 69306
rect 90014 69144 92514 69306
rect 92682 69144 95090 69306
rect 95258 69144 97666 69306
rect 97834 69144 100334 69306
rect 100502 69144 102910 69306
rect 103078 69144 105486 69306
rect 105654 69144 108154 69306
rect 108322 69144 110730 69306
rect 110898 69144 113306 69306
rect 113474 69144 115974 69306
rect 116142 69144 118550 69306
rect 118718 69144 119396 69306
rect 572 856 119396 69144
rect 682 2 1618 856
rect 1786 2 2814 856
rect 2982 2 4010 856
rect 4178 2 5206 856
rect 5374 2 6310 856
rect 6478 2 7506 856
rect 7674 2 8702 856
rect 8870 2 9898 856
rect 10066 2 11094 856
rect 11262 2 12198 856
rect 12366 2 13394 856
rect 13562 2 14590 856
rect 14758 2 15786 856
rect 15954 2 16890 856
rect 17058 2 18086 856
rect 18254 2 19282 856
rect 19450 2 20478 856
rect 20646 2 21674 856
rect 21842 2 22778 856
rect 22946 2 23974 856
rect 24142 2 25170 856
rect 25338 2 26366 856
rect 26534 2 27562 856
rect 27730 2 28666 856
rect 28834 2 29862 856
rect 30030 2 31058 856
rect 31226 2 32254 856
rect 32422 2 33358 856
rect 33526 2 34554 856
rect 34722 2 35750 856
rect 35918 2 36946 856
rect 37114 2 38142 856
rect 38310 2 39246 856
rect 39414 2 40442 856
rect 40610 2 41638 856
rect 41806 2 42834 856
rect 43002 2 44030 856
rect 44198 2 45134 856
rect 45302 2 46330 856
rect 46498 2 47526 856
rect 47694 2 48722 856
rect 48890 2 49826 856
rect 49994 2 51022 856
rect 51190 2 52218 856
rect 52386 2 53414 856
rect 53582 2 54610 856
rect 54778 2 55714 856
rect 55882 2 56910 856
rect 57078 2 58106 856
rect 58274 2 59302 856
rect 59470 2 60498 856
rect 60666 2 61602 856
rect 61770 2 62798 856
rect 62966 2 63994 856
rect 64162 2 65190 856
rect 65358 2 66294 856
rect 66462 2 67490 856
rect 67658 2 68686 856
rect 68854 2 69882 856
rect 70050 2 71078 856
rect 71246 2 72182 856
rect 72350 2 73378 856
rect 73546 2 74574 856
rect 74742 2 75770 856
rect 75938 2 76874 856
rect 77042 2 78070 856
rect 78238 2 79266 856
rect 79434 2 80462 856
rect 80630 2 81658 856
rect 81826 2 82762 856
rect 82930 2 83958 856
rect 84126 2 85154 856
rect 85322 2 86350 856
rect 86518 2 87546 856
rect 87714 2 88650 856
rect 88818 2 89846 856
rect 90014 2 91042 856
rect 91210 2 92238 856
rect 92406 2 93342 856
rect 93510 2 94538 856
rect 94706 2 95734 856
rect 95902 2 96930 856
rect 97098 2 98126 856
rect 98294 2 99230 856
rect 99398 2 100426 856
rect 100594 2 101622 856
rect 101790 2 102818 856
rect 102986 2 104014 856
rect 104182 2 105118 856
rect 105286 2 106314 856
rect 106482 2 107510 856
rect 107678 2 108706 856
rect 108874 2 109810 856
rect 109978 2 111006 856
rect 111174 2 112202 856
rect 112370 2 113398 856
rect 113566 2 114594 856
rect 114762 2 115698 856
rect 115866 2 116894 856
rect 117062 2 118090 856
rect 118258 2 119286 856
<< metal3 >>
rect 0 69096 800 69216
rect 0 67464 800 67584
rect 0 65832 800 65952
rect 0 64200 800 64320
rect 0 62568 800 62688
rect 0 60936 800 61056
rect 0 59304 800 59424
rect 0 57672 800 57792
rect 0 56040 800 56160
rect 0 54408 800 54528
rect 0 52776 800 52896
rect 0 51144 800 51264
rect 0 49512 800 49632
rect 0 47880 800 48000
rect 0 46248 800 46368
rect 0 44616 800 44736
rect 0 42984 800 43104
rect 0 41352 800 41472
rect 0 39720 800 39840
rect 0 38088 800 38208
rect 0 36456 800 36576
rect 0 34824 800 34944
rect 0 33192 800 33312
rect 0 31560 800 31680
rect 0 29928 800 30048
rect 0 28296 800 28416
rect 0 26664 800 26784
rect 0 25032 800 25152
rect 0 23400 800 23520
rect 0 21768 800 21888
rect 0 20136 800 20256
rect 0 18504 800 18624
rect 0 16872 800 16992
rect 0 15240 800 15360
rect 0 13608 800 13728
rect 0 11976 800 12096
rect 0 10344 800 10464
rect 0 8712 800 8832
rect 0 7080 800 7200
rect 0 5448 800 5568
rect 0 3816 800 3936
rect 0 2184 800 2304
rect 0 688 800 808
<< obsm3 >>
rect 880 69016 116183 69189
rect 800 67664 116183 69016
rect 880 67384 116183 67664
rect 800 66032 116183 67384
rect 880 65752 116183 66032
rect 800 64400 116183 65752
rect 880 64120 116183 64400
rect 800 62768 116183 64120
rect 880 62488 116183 62768
rect 800 61136 116183 62488
rect 880 60856 116183 61136
rect 800 59504 116183 60856
rect 880 59224 116183 59504
rect 800 57872 116183 59224
rect 880 57592 116183 57872
rect 800 56240 116183 57592
rect 880 55960 116183 56240
rect 800 54608 116183 55960
rect 880 54328 116183 54608
rect 800 52976 116183 54328
rect 880 52696 116183 52976
rect 800 51344 116183 52696
rect 880 51064 116183 51344
rect 800 49712 116183 51064
rect 880 49432 116183 49712
rect 800 48080 116183 49432
rect 880 47800 116183 48080
rect 800 46448 116183 47800
rect 880 46168 116183 46448
rect 800 44816 116183 46168
rect 880 44536 116183 44816
rect 800 43184 116183 44536
rect 880 42904 116183 43184
rect 800 41552 116183 42904
rect 880 41272 116183 41552
rect 800 39920 116183 41272
rect 880 39640 116183 39920
rect 800 38288 116183 39640
rect 880 38008 116183 38288
rect 800 36656 116183 38008
rect 880 36376 116183 36656
rect 800 35024 116183 36376
rect 880 34744 116183 35024
rect 800 33392 116183 34744
rect 880 33112 116183 33392
rect 800 31760 116183 33112
rect 880 31480 116183 31760
rect 800 30128 116183 31480
rect 880 29848 116183 30128
rect 800 28496 116183 29848
rect 880 28216 116183 28496
rect 800 26864 116183 28216
rect 880 26584 116183 26864
rect 800 25232 116183 26584
rect 880 24952 116183 25232
rect 800 23600 116183 24952
rect 880 23320 116183 23600
rect 800 21968 116183 23320
rect 880 21688 116183 21968
rect 800 20336 116183 21688
rect 880 20056 116183 20336
rect 800 18704 116183 20056
rect 880 18424 116183 18704
rect 800 17072 116183 18424
rect 880 16792 116183 17072
rect 800 15440 116183 16792
rect 880 15160 116183 15440
rect 800 13808 116183 15160
rect 880 13528 116183 13808
rect 800 12176 116183 13528
rect 880 11896 116183 12176
rect 800 10544 116183 11896
rect 880 10264 116183 10544
rect 800 8912 116183 10264
rect 880 8632 116183 8912
rect 800 7280 116183 8632
rect 880 7000 116183 7280
rect 800 5648 116183 7000
rect 880 5368 116183 5648
rect 800 4016 116183 5368
rect 880 3736 116183 4016
rect 800 2384 116183 3736
rect 880 2104 116183 2384
rect 800 888 116183 2104
rect 880 715 116183 888
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
rect 81008 2128 81328 67504
rect 96368 2128 96688 67504
rect 111728 2128 112048 67504
<< obsm4 >>
rect 19379 4523 19488 67285
rect 19968 4523 34848 67285
rect 35328 4523 50208 67285
rect 50688 4523 65568 67285
rect 66048 4523 80928 67285
rect 81408 4523 96288 67285
rect 96768 4523 103349 67285
<< labels >>
rlabel metal3 s 0 2184 800 2304 6 addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 addr1[9]
port 10 nsew signal output
rlabel metal3 s 0 688 800 808 6 csb1
port 11 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 dout1[0]
port 12 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 dout1[10]
port 13 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 dout1[11]
port 14 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 dout1[12]
port 15 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 dout1[13]
port 16 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 dout1[14]
port 17 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 dout1[15]
port 18 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 dout1[16]
port 19 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 dout1[17]
port 20 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 dout1[18]
port 21 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 dout1[19]
port 22 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 dout1[1]
port 23 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 dout1[20]
port 24 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 dout1[21]
port 25 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 dout1[22]
port 26 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 dout1[23]
port 27 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 dout1[24]
port 28 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 dout1[25]
port 29 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 dout1[26]
port 30 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 dout1[27]
port 31 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 dout1[28]
port 32 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 dout1[29]
port 33 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 dout1[2]
port 34 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 dout1[30]
port 35 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 dout1[31]
port 36 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 dout1[3]
port 37 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 dout1[4]
port 38 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 dout1[5]
port 39 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 dout1[6]
port 40 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 dout1[7]
port 41 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 dout1[8]
port 42 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 dout1[9]
port 43 nsew signal input
rlabel metal2 s 92570 69200 92626 70000 6 io_oeb[0]
port 44 nsew signal output
rlabel metal2 s 118606 69200 118662 70000 6 io_oeb[10]
port 45 nsew signal output
rlabel metal2 s 95146 69200 95202 70000 6 io_oeb[1]
port 46 nsew signal output
rlabel metal2 s 97722 69200 97778 70000 6 io_oeb[2]
port 47 nsew signal output
rlabel metal2 s 100390 69200 100446 70000 6 io_oeb[3]
port 48 nsew signal output
rlabel metal2 s 102966 69200 103022 70000 6 io_oeb[4]
port 49 nsew signal output
rlabel metal2 s 105542 69200 105598 70000 6 io_oeb[5]
port 50 nsew signal output
rlabel metal2 s 108210 69200 108266 70000 6 io_oeb[6]
port 51 nsew signal output
rlabel metal2 s 110786 69200 110842 70000 6 io_oeb[7]
port 52 nsew signal output
rlabel metal2 s 113362 69200 113418 70000 6 io_oeb[8]
port 53 nsew signal output
rlabel metal2 s 116030 69200 116086 70000 6 io_oeb[9]
port 54 nsew signal output
rlabel metal2 s 570 0 626 800 6 io_wbs_ack
port 55 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 io_wbs_adr[0]
port 56 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 io_wbs_adr[10]
port 57 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 io_wbs_adr[11]
port 58 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 io_wbs_adr[12]
port 59 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 io_wbs_adr[13]
port 60 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 io_wbs_adr[14]
port 61 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 io_wbs_adr[15]
port 62 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 io_wbs_adr[16]
port 63 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 io_wbs_adr[17]
port 64 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 io_wbs_adr[18]
port 65 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 io_wbs_adr[19]
port 66 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 io_wbs_adr[1]
port 67 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 io_wbs_adr[20]
port 68 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 io_wbs_adr[21]
port 69 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 io_wbs_adr[22]
port 70 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 io_wbs_adr[23]
port 71 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 io_wbs_adr[24]
port 72 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 io_wbs_adr[25]
port 73 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 io_wbs_adr[26]
port 74 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 io_wbs_adr[27]
port 75 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 io_wbs_adr[28]
port 76 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 io_wbs_adr[29]
port 77 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 io_wbs_adr[2]
port 78 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 io_wbs_adr[30]
port 79 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 io_wbs_adr[31]
port 80 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 io_wbs_adr[3]
port 81 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 io_wbs_adr[4]
port 82 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 io_wbs_adr[5]
port 83 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 io_wbs_adr[6]
port 84 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 io_wbs_adr[7]
port 85 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 io_wbs_adr[8]
port 86 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 io_wbs_adr[9]
port 87 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 io_wbs_clk
port 88 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 io_wbs_cyc
port 89 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 io_wbs_datrd[0]
port 90 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 io_wbs_datrd[10]
port 91 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 io_wbs_datrd[11]
port 92 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 io_wbs_datrd[12]
port 93 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 io_wbs_datrd[13]
port 94 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 io_wbs_datrd[14]
port 95 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 io_wbs_datrd[15]
port 96 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 io_wbs_datrd[16]
port 97 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 io_wbs_datrd[17]
port 98 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 io_wbs_datrd[18]
port 99 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 io_wbs_datrd[19]
port 100 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 io_wbs_datrd[1]
port 101 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 io_wbs_datrd[20]
port 102 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 io_wbs_datrd[21]
port 103 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 io_wbs_datrd[22]
port 104 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 io_wbs_datrd[23]
port 105 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 io_wbs_datrd[24]
port 106 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 io_wbs_datrd[25]
port 107 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 io_wbs_datrd[26]
port 108 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 io_wbs_datrd[27]
port 109 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 io_wbs_datrd[28]
port 110 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 io_wbs_datrd[29]
port 111 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 io_wbs_datrd[2]
port 112 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 io_wbs_datrd[30]
port 113 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 io_wbs_datrd[31]
port 114 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_wbs_datrd[3]
port 115 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 io_wbs_datrd[4]
port 116 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 io_wbs_datrd[5]
port 117 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_wbs_datrd[6]
port 118 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 io_wbs_datrd[7]
port 119 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 io_wbs_datrd[8]
port 120 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 io_wbs_datrd[9]
port 121 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 io_wbs_datwr[0]
port 122 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 io_wbs_datwr[10]
port 123 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 io_wbs_datwr[11]
port 124 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 io_wbs_datwr[12]
port 125 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 io_wbs_datwr[13]
port 126 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 io_wbs_datwr[14]
port 127 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 io_wbs_datwr[15]
port 128 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 io_wbs_datwr[16]
port 129 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 io_wbs_datwr[17]
port 130 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 io_wbs_datwr[18]
port 131 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 io_wbs_datwr[19]
port 132 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 io_wbs_datwr[1]
port 133 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 io_wbs_datwr[20]
port 134 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 io_wbs_datwr[21]
port 135 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 io_wbs_datwr[22]
port 136 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 io_wbs_datwr[23]
port 137 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 io_wbs_datwr[24]
port 138 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 io_wbs_datwr[25]
port 139 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 io_wbs_datwr[26]
port 140 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 io_wbs_datwr[27]
port 141 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 io_wbs_datwr[28]
port 142 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 io_wbs_datwr[29]
port 143 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 io_wbs_datwr[2]
port 144 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 io_wbs_datwr[30]
port 145 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 io_wbs_datwr[31]
port 146 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 io_wbs_datwr[3]
port 147 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 io_wbs_datwr[4]
port 148 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 io_wbs_datwr[5]
port 149 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 io_wbs_datwr[6]
port 150 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 io_wbs_datwr[7]
port 151 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 io_wbs_datwr[8]
port 152 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 io_wbs_datwr[9]
port 153 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 io_wbs_rst
port 154 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 io_wbs_stb
port 155 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 io_wbs_we
port 156 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 157 nsew power input
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 157 nsew power input
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 157 nsew power input
rlabel metal4 s 96368 2128 96688 67504 6 vccd1
port 157 nsew power input
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 158 nsew ground input
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 158 nsew ground input
rlabel metal4 s 81008 2128 81328 67504 6 vssd1
port 158 nsew ground input
rlabel metal4 s 111728 2128 112048 67504 6 vssd1
port 158 nsew ground input
rlabel metal2 s 9126 69200 9182 70000 6 wfg_drive_pat_dout_o[0]
port 159 nsew signal output
rlabel metal2 s 35162 69200 35218 70000 6 wfg_drive_pat_dout_o[10]
port 160 nsew signal output
rlabel metal2 s 37738 69200 37794 70000 6 wfg_drive_pat_dout_o[11]
port 161 nsew signal output
rlabel metal2 s 40406 69200 40462 70000 6 wfg_drive_pat_dout_o[12]
port 162 nsew signal output
rlabel metal2 s 42982 69200 43038 70000 6 wfg_drive_pat_dout_o[13]
port 163 nsew signal output
rlabel metal2 s 45558 69200 45614 70000 6 wfg_drive_pat_dout_o[14]
port 164 nsew signal output
rlabel metal2 s 48226 69200 48282 70000 6 wfg_drive_pat_dout_o[15]
port 165 nsew signal output
rlabel metal2 s 50802 69200 50858 70000 6 wfg_drive_pat_dout_o[16]
port 166 nsew signal output
rlabel metal2 s 53378 69200 53434 70000 6 wfg_drive_pat_dout_o[17]
port 167 nsew signal output
rlabel metal2 s 56046 69200 56102 70000 6 wfg_drive_pat_dout_o[18]
port 168 nsew signal output
rlabel metal2 s 58622 69200 58678 70000 6 wfg_drive_pat_dout_o[19]
port 169 nsew signal output
rlabel metal2 s 11702 69200 11758 70000 6 wfg_drive_pat_dout_o[1]
port 170 nsew signal output
rlabel metal2 s 61290 69200 61346 70000 6 wfg_drive_pat_dout_o[20]
port 171 nsew signal output
rlabel metal2 s 63866 69200 63922 70000 6 wfg_drive_pat_dout_o[21]
port 172 nsew signal output
rlabel metal2 s 66442 69200 66498 70000 6 wfg_drive_pat_dout_o[22]
port 173 nsew signal output
rlabel metal2 s 69110 69200 69166 70000 6 wfg_drive_pat_dout_o[23]
port 174 nsew signal output
rlabel metal2 s 71686 69200 71742 70000 6 wfg_drive_pat_dout_o[24]
port 175 nsew signal output
rlabel metal2 s 74262 69200 74318 70000 6 wfg_drive_pat_dout_o[25]
port 176 nsew signal output
rlabel metal2 s 76930 69200 76986 70000 6 wfg_drive_pat_dout_o[26]
port 177 nsew signal output
rlabel metal2 s 79506 69200 79562 70000 6 wfg_drive_pat_dout_o[27]
port 178 nsew signal output
rlabel metal2 s 82082 69200 82138 70000 6 wfg_drive_pat_dout_o[28]
port 179 nsew signal output
rlabel metal2 s 84750 69200 84806 70000 6 wfg_drive_pat_dout_o[29]
port 180 nsew signal output
rlabel metal2 s 14278 69200 14334 70000 6 wfg_drive_pat_dout_o[2]
port 181 nsew signal output
rlabel metal2 s 87326 69200 87382 70000 6 wfg_drive_pat_dout_o[30]
port 182 nsew signal output
rlabel metal2 s 89902 69200 89958 70000 6 wfg_drive_pat_dout_o[31]
port 183 nsew signal output
rlabel metal2 s 16946 69200 17002 70000 6 wfg_drive_pat_dout_o[3]
port 184 nsew signal output
rlabel metal2 s 19522 69200 19578 70000 6 wfg_drive_pat_dout_o[4]
port 185 nsew signal output
rlabel metal2 s 22098 69200 22154 70000 6 wfg_drive_pat_dout_o[5]
port 186 nsew signal output
rlabel metal2 s 24766 69200 24822 70000 6 wfg_drive_pat_dout_o[6]
port 187 nsew signal output
rlabel metal2 s 27342 69200 27398 70000 6 wfg_drive_pat_dout_o[7]
port 188 nsew signal output
rlabel metal2 s 29918 69200 29974 70000 6 wfg_drive_pat_dout_o[8]
port 189 nsew signal output
rlabel metal2 s 32586 69200 32642 70000 6 wfg_drive_pat_dout_o[9]
port 190 nsew signal output
rlabel metal2 s 1306 69200 1362 70000 6 wfg_drive_spi_cs_no
port 191 nsew signal output
rlabel metal2 s 3882 69200 3938 70000 6 wfg_drive_spi_sclk_o
port 192 nsew signal output
rlabel metal2 s 6458 69200 6514 70000 6 wfg_drive_spi_sdo_o
port 193 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23342254
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/user_proj_wfg/runs/user_proj_wfg/results/finishing/wfg_top.magic.gds
string GDS_START 1362936
<< end >>

