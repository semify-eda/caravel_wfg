magic
tech sky130A
magscale 1 2
timestamp 1657112955
<< obsli1 >>
rect 1104 2159 148856 107729
<< obsm1 >>
rect 658 1640 149210 107760
<< metal2 >>
rect 1582 109200 1638 110000
rect 4802 109200 4858 110000
rect 8022 109200 8078 110000
rect 11334 109200 11390 110000
rect 14554 109200 14610 110000
rect 17866 109200 17922 110000
rect 21086 109200 21142 110000
rect 24398 109200 24454 110000
rect 27618 109200 27674 110000
rect 30838 109200 30894 110000
rect 34150 109200 34206 110000
rect 37370 109200 37426 110000
rect 40682 109200 40738 110000
rect 43902 109200 43958 110000
rect 47214 109200 47270 110000
rect 50434 109200 50490 110000
rect 53654 109200 53710 110000
rect 56966 109200 57022 110000
rect 60186 109200 60242 110000
rect 63498 109200 63554 110000
rect 66718 109200 66774 110000
rect 70030 109200 70086 110000
rect 73250 109200 73306 110000
rect 76562 109200 76618 110000
rect 79782 109200 79838 110000
rect 83002 109200 83058 110000
rect 86314 109200 86370 110000
rect 89534 109200 89590 110000
rect 92846 109200 92902 110000
rect 96066 109200 96122 110000
rect 99378 109200 99434 110000
rect 102598 109200 102654 110000
rect 105818 109200 105874 110000
rect 109130 109200 109186 110000
rect 112350 109200 112406 110000
rect 115662 109200 115718 110000
rect 118882 109200 118938 110000
rect 122194 109200 122250 110000
rect 125414 109200 125470 110000
rect 128634 109200 128690 110000
rect 131946 109200 132002 110000
rect 135166 109200 135222 110000
rect 138478 109200 138534 110000
rect 141698 109200 141754 110000
rect 145010 109200 145066 110000
rect 148230 109200 148286 110000
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4986 0 5042 800
rect 6458 0 6514 800
rect 7930 0 7986 800
rect 9402 0 9458 800
rect 10874 0 10930 800
rect 12346 0 12402 800
rect 13818 0 13874 800
rect 15290 0 15346 800
rect 16762 0 16818 800
rect 18234 0 18290 800
rect 19706 0 19762 800
rect 21178 0 21234 800
rect 22650 0 22706 800
rect 24122 0 24178 800
rect 25594 0 25650 800
rect 27066 0 27122 800
rect 28538 0 28594 800
rect 30010 0 30066 800
rect 31482 0 31538 800
rect 32954 0 33010 800
rect 34426 0 34482 800
rect 35898 0 35954 800
rect 37370 0 37426 800
rect 38842 0 38898 800
rect 40314 0 40370 800
rect 41786 0 41842 800
rect 43258 0 43314 800
rect 44730 0 44786 800
rect 46202 0 46258 800
rect 47674 0 47730 800
rect 49146 0 49202 800
rect 50618 0 50674 800
rect 52090 0 52146 800
rect 53562 0 53618 800
rect 55034 0 55090 800
rect 56506 0 56562 800
rect 57978 0 58034 800
rect 59450 0 59506 800
rect 60922 0 60978 800
rect 62394 0 62450 800
rect 63866 0 63922 800
rect 65338 0 65394 800
rect 66810 0 66866 800
rect 68282 0 68338 800
rect 69754 0 69810 800
rect 71226 0 71282 800
rect 72698 0 72754 800
rect 74170 0 74226 800
rect 75642 0 75698 800
rect 77022 0 77078 800
rect 78494 0 78550 800
rect 79966 0 80022 800
rect 81438 0 81494 800
rect 82910 0 82966 800
rect 84382 0 84438 800
rect 85854 0 85910 800
rect 87326 0 87382 800
rect 88798 0 88854 800
rect 90270 0 90326 800
rect 91742 0 91798 800
rect 93214 0 93270 800
rect 94686 0 94742 800
rect 96158 0 96214 800
rect 97630 0 97686 800
rect 99102 0 99158 800
rect 100574 0 100630 800
rect 102046 0 102102 800
rect 103518 0 103574 800
rect 104990 0 105046 800
rect 106462 0 106518 800
rect 107934 0 107990 800
rect 109406 0 109462 800
rect 110878 0 110934 800
rect 112350 0 112406 800
rect 113822 0 113878 800
rect 115294 0 115350 800
rect 116766 0 116822 800
rect 118238 0 118294 800
rect 119710 0 119766 800
rect 121182 0 121238 800
rect 122654 0 122710 800
rect 124126 0 124182 800
rect 125598 0 125654 800
rect 127070 0 127126 800
rect 128542 0 128598 800
rect 130014 0 130070 800
rect 131486 0 131542 800
rect 132958 0 133014 800
rect 134430 0 134486 800
rect 135902 0 135958 800
rect 137374 0 137430 800
rect 138846 0 138902 800
rect 140318 0 140374 800
rect 141790 0 141846 800
rect 143262 0 143318 800
rect 144734 0 144790 800
rect 146206 0 146262 800
rect 147678 0 147734 800
rect 149150 0 149206 800
<< obsm2 >>
rect 664 109144 1526 109200
rect 1694 109144 4746 109200
rect 4914 109144 7966 109200
rect 8134 109144 11278 109200
rect 11446 109144 14498 109200
rect 14666 109144 17810 109200
rect 17978 109144 21030 109200
rect 21198 109144 24342 109200
rect 24510 109144 27562 109200
rect 27730 109144 30782 109200
rect 30950 109144 34094 109200
rect 34262 109144 37314 109200
rect 37482 109144 40626 109200
rect 40794 109144 43846 109200
rect 44014 109144 47158 109200
rect 47326 109144 50378 109200
rect 50546 109144 53598 109200
rect 53766 109144 56910 109200
rect 57078 109144 60130 109200
rect 60298 109144 63442 109200
rect 63610 109144 66662 109200
rect 66830 109144 69974 109200
rect 70142 109144 73194 109200
rect 73362 109144 76506 109200
rect 76674 109144 79726 109200
rect 79894 109144 82946 109200
rect 83114 109144 86258 109200
rect 86426 109144 89478 109200
rect 89646 109144 92790 109200
rect 92958 109144 96010 109200
rect 96178 109144 99322 109200
rect 99490 109144 102542 109200
rect 102710 109144 105762 109200
rect 105930 109144 109074 109200
rect 109242 109144 112294 109200
rect 112462 109144 115606 109200
rect 115774 109144 118826 109200
rect 118994 109144 122138 109200
rect 122306 109144 125358 109200
rect 125526 109144 128578 109200
rect 128746 109144 131890 109200
rect 132058 109144 135110 109200
rect 135278 109144 138422 109200
rect 138590 109144 141642 109200
rect 141810 109144 144954 109200
rect 145122 109144 148174 109200
rect 148342 109144 149204 109200
rect 664 856 149204 109144
rect 774 734 1986 856
rect 2154 734 3458 856
rect 3626 734 4930 856
rect 5098 734 6402 856
rect 6570 734 7874 856
rect 8042 734 9346 856
rect 9514 734 10818 856
rect 10986 734 12290 856
rect 12458 734 13762 856
rect 13930 734 15234 856
rect 15402 734 16706 856
rect 16874 734 18178 856
rect 18346 734 19650 856
rect 19818 734 21122 856
rect 21290 734 22594 856
rect 22762 734 24066 856
rect 24234 734 25538 856
rect 25706 734 27010 856
rect 27178 734 28482 856
rect 28650 734 29954 856
rect 30122 734 31426 856
rect 31594 734 32898 856
rect 33066 734 34370 856
rect 34538 734 35842 856
rect 36010 734 37314 856
rect 37482 734 38786 856
rect 38954 734 40258 856
rect 40426 734 41730 856
rect 41898 734 43202 856
rect 43370 734 44674 856
rect 44842 734 46146 856
rect 46314 734 47618 856
rect 47786 734 49090 856
rect 49258 734 50562 856
rect 50730 734 52034 856
rect 52202 734 53506 856
rect 53674 734 54978 856
rect 55146 734 56450 856
rect 56618 734 57922 856
rect 58090 734 59394 856
rect 59562 734 60866 856
rect 61034 734 62338 856
rect 62506 734 63810 856
rect 63978 734 65282 856
rect 65450 734 66754 856
rect 66922 734 68226 856
rect 68394 734 69698 856
rect 69866 734 71170 856
rect 71338 734 72642 856
rect 72810 734 74114 856
rect 74282 734 75586 856
rect 75754 734 76966 856
rect 77134 734 78438 856
rect 78606 734 79910 856
rect 80078 734 81382 856
rect 81550 734 82854 856
rect 83022 734 84326 856
rect 84494 734 85798 856
rect 85966 734 87270 856
rect 87438 734 88742 856
rect 88910 734 90214 856
rect 90382 734 91686 856
rect 91854 734 93158 856
rect 93326 734 94630 856
rect 94798 734 96102 856
rect 96270 734 97574 856
rect 97742 734 99046 856
rect 99214 734 100518 856
rect 100686 734 101990 856
rect 102158 734 103462 856
rect 103630 734 104934 856
rect 105102 734 106406 856
rect 106574 734 107878 856
rect 108046 734 109350 856
rect 109518 734 110822 856
rect 110990 734 112294 856
rect 112462 734 113766 856
rect 113934 734 115238 856
rect 115406 734 116710 856
rect 116878 734 118182 856
rect 118350 734 119654 856
rect 119822 734 121126 856
rect 121294 734 122598 856
rect 122766 734 124070 856
rect 124238 734 125542 856
rect 125710 734 127014 856
rect 127182 734 128486 856
rect 128654 734 129958 856
rect 130126 734 131430 856
rect 131598 734 132902 856
rect 133070 734 134374 856
rect 134542 734 135846 856
rect 136014 734 137318 856
rect 137486 734 138790 856
rect 138958 734 140262 856
rect 140430 734 141734 856
rect 141902 734 143206 856
rect 143374 734 144678 856
rect 144846 734 146150 856
rect 146318 734 147622 856
rect 147790 734 149094 856
<< metal3 >>
rect 0 108672 800 108792
rect 0 106088 800 106208
rect 0 103504 800 103624
rect 0 100920 800 101040
rect 0 98336 800 98456
rect 0 95888 800 96008
rect 0 93304 800 93424
rect 0 90720 800 90840
rect 0 88136 800 88256
rect 0 85552 800 85672
rect 0 83104 800 83224
rect 0 80520 800 80640
rect 0 77936 800 78056
rect 0 75352 800 75472
rect 0 72768 800 72888
rect 0 70184 800 70304
rect 0 67736 800 67856
rect 0 65152 800 65272
rect 0 62568 800 62688
rect 0 59984 800 60104
rect 0 57400 800 57520
rect 0 54952 800 55072
rect 0 52368 800 52488
rect 0 49784 800 49904
rect 0 47200 800 47320
rect 0 44616 800 44736
rect 0 42168 800 42288
rect 0 39584 800 39704
rect 0 37000 800 37120
rect 0 34416 800 34536
rect 0 31832 800 31952
rect 0 29248 800 29368
rect 0 26800 800 26920
rect 0 24216 800 24336
rect 0 21632 800 21752
rect 0 19048 800 19168
rect 0 16464 800 16584
rect 0 14016 800 14136
rect 0 11432 800 11552
rect 0 8848 800 8968
rect 0 6264 800 6384
rect 0 3680 800 3800
rect 0 1232 800 1352
<< obsm3 >>
rect 880 108592 146543 108765
rect 800 106288 146543 108592
rect 880 106008 146543 106288
rect 800 103704 146543 106008
rect 880 103424 146543 103704
rect 800 101120 146543 103424
rect 880 100840 146543 101120
rect 800 98536 146543 100840
rect 880 98256 146543 98536
rect 800 96088 146543 98256
rect 880 95808 146543 96088
rect 800 93504 146543 95808
rect 880 93224 146543 93504
rect 800 90920 146543 93224
rect 880 90640 146543 90920
rect 800 88336 146543 90640
rect 880 88056 146543 88336
rect 800 85752 146543 88056
rect 880 85472 146543 85752
rect 800 83304 146543 85472
rect 880 83024 146543 83304
rect 800 80720 146543 83024
rect 880 80440 146543 80720
rect 800 78136 146543 80440
rect 880 77856 146543 78136
rect 800 75552 146543 77856
rect 880 75272 146543 75552
rect 800 72968 146543 75272
rect 880 72688 146543 72968
rect 800 70384 146543 72688
rect 880 70104 146543 70384
rect 800 67936 146543 70104
rect 880 67656 146543 67936
rect 800 65352 146543 67656
rect 880 65072 146543 65352
rect 800 62768 146543 65072
rect 880 62488 146543 62768
rect 800 60184 146543 62488
rect 880 59904 146543 60184
rect 800 57600 146543 59904
rect 880 57320 146543 57600
rect 800 55152 146543 57320
rect 880 54872 146543 55152
rect 800 52568 146543 54872
rect 880 52288 146543 52568
rect 800 49984 146543 52288
rect 880 49704 146543 49984
rect 800 47400 146543 49704
rect 880 47120 146543 47400
rect 800 44816 146543 47120
rect 880 44536 146543 44816
rect 800 42368 146543 44536
rect 880 42088 146543 42368
rect 800 39784 146543 42088
rect 880 39504 146543 39784
rect 800 37200 146543 39504
rect 880 36920 146543 37200
rect 800 34616 146543 36920
rect 880 34336 146543 34616
rect 800 32032 146543 34336
rect 880 31752 146543 32032
rect 800 29448 146543 31752
rect 880 29168 146543 29448
rect 800 27000 146543 29168
rect 880 26720 146543 27000
rect 800 24416 146543 26720
rect 880 24136 146543 24416
rect 800 21832 146543 24136
rect 880 21552 146543 21832
rect 800 19248 146543 21552
rect 880 18968 146543 19248
rect 800 16664 146543 18968
rect 880 16384 146543 16664
rect 800 14216 146543 16384
rect 880 13936 146543 14216
rect 800 11632 146543 13936
rect 880 11352 146543 11632
rect 800 9048 146543 11352
rect 880 8768 146543 9048
rect 800 6464 146543 8768
rect 880 6184 146543 6464
rect 800 3880 146543 6184
rect 880 3600 146543 3880
rect 800 1432 146543 3600
rect 880 1259 146543 1432
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
rect 111728 2128 112048 107760
rect 127088 2128 127408 107760
rect 142448 2128 142768 107760
<< obsm4 >>
rect 5763 2891 19488 107405
rect 19968 2891 34848 107405
rect 35328 2891 50208 107405
rect 50688 2891 65568 107405
rect 66048 2891 80928 107405
rect 81408 2891 96288 107405
rect 96768 2891 111648 107405
rect 112128 2891 127008 107405
rect 127488 2891 129477 107405
<< labels >>
rlabel metal3 s 0 3680 800 3800 6 addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 addr1[9]
port 10 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 csb1
port 11 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 dout1[0]
port 12 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 dout1[10]
port 13 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 dout1[11]
port 14 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 dout1[12]
port 15 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 dout1[13]
port 16 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 dout1[14]
port 17 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 dout1[15]
port 18 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 dout1[16]
port 19 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 dout1[17]
port 20 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 dout1[18]
port 21 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 dout1[19]
port 22 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 dout1[1]
port 23 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 dout1[20]
port 24 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 dout1[21]
port 25 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 dout1[22]
port 26 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 dout1[23]
port 27 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 dout1[24]
port 28 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 dout1[25]
port 29 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 dout1[26]
port 30 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 dout1[27]
port 31 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 dout1[28]
port 32 nsew signal input
rlabel metal3 s 0 103504 800 103624 6 dout1[29]
port 33 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 dout1[2]
port 34 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 dout1[30]
port 35 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 dout1[31]
port 36 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 dout1[3]
port 37 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 dout1[4]
port 38 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 dout1[5]
port 39 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 dout1[6]
port 40 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 dout1[7]
port 41 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 dout1[8]
port 42 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 dout1[9]
port 43 nsew signal input
rlabel metal2 s 115662 109200 115718 110000 6 io_oeb[0]
port 44 nsew signal output
rlabel metal2 s 148230 109200 148286 110000 6 io_oeb[10]
port 45 nsew signal output
rlabel metal2 s 118882 109200 118938 110000 6 io_oeb[1]
port 46 nsew signal output
rlabel metal2 s 122194 109200 122250 110000 6 io_oeb[2]
port 47 nsew signal output
rlabel metal2 s 125414 109200 125470 110000 6 io_oeb[3]
port 48 nsew signal output
rlabel metal2 s 128634 109200 128690 110000 6 io_oeb[4]
port 49 nsew signal output
rlabel metal2 s 131946 109200 132002 110000 6 io_oeb[5]
port 50 nsew signal output
rlabel metal2 s 135166 109200 135222 110000 6 io_oeb[6]
port 51 nsew signal output
rlabel metal2 s 138478 109200 138534 110000 6 io_oeb[7]
port 52 nsew signal output
rlabel metal2 s 141698 109200 141754 110000 6 io_oeb[8]
port 53 nsew signal output
rlabel metal2 s 145010 109200 145066 110000 6 io_oeb[9]
port 54 nsew signal output
rlabel metal2 s 662 0 718 800 6 io_wbs_ack
port 55 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 io_wbs_adr[0]
port 56 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 io_wbs_adr[10]
port 57 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 io_wbs_adr[11]
port 58 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 io_wbs_adr[12]
port 59 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 io_wbs_adr[13]
port 60 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 io_wbs_adr[14]
port 61 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 io_wbs_adr[15]
port 62 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 io_wbs_adr[16]
port 63 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 io_wbs_adr[17]
port 64 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 io_wbs_adr[18]
port 65 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 io_wbs_adr[19]
port 66 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 io_wbs_adr[1]
port 67 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 io_wbs_adr[20]
port 68 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 io_wbs_adr[21]
port 69 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 io_wbs_adr[22]
port 70 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 io_wbs_adr[23]
port 71 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 io_wbs_adr[24]
port 72 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 io_wbs_adr[25]
port 73 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 io_wbs_adr[26]
port 74 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 io_wbs_adr[27]
port 75 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 io_wbs_adr[28]
port 76 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 io_wbs_adr[29]
port 77 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 io_wbs_adr[2]
port 78 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 io_wbs_adr[30]
port 79 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 io_wbs_adr[31]
port 80 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 io_wbs_adr[3]
port 81 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 io_wbs_adr[4]
port 82 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 io_wbs_adr[5]
port 83 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 io_wbs_adr[6]
port 84 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 io_wbs_adr[7]
port 85 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 io_wbs_adr[8]
port 86 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 io_wbs_adr[9]
port 87 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 io_wbs_clk
port 88 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 io_wbs_cyc
port 89 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_wbs_datrd[0]
port 90 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 io_wbs_datrd[10]
port 91 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 io_wbs_datrd[11]
port 92 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 io_wbs_datrd[12]
port 93 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 io_wbs_datrd[13]
port 94 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 io_wbs_datrd[14]
port 95 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 io_wbs_datrd[15]
port 96 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 io_wbs_datrd[16]
port 97 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 io_wbs_datrd[17]
port 98 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 io_wbs_datrd[18]
port 99 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 io_wbs_datrd[19]
port 100 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 io_wbs_datrd[1]
port 101 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 io_wbs_datrd[20]
port 102 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 io_wbs_datrd[21]
port 103 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 io_wbs_datrd[22]
port 104 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 io_wbs_datrd[23]
port 105 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 io_wbs_datrd[24]
port 106 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 io_wbs_datrd[25]
port 107 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 io_wbs_datrd[26]
port 108 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 io_wbs_datrd[27]
port 109 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 io_wbs_datrd[28]
port 110 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 io_wbs_datrd[29]
port 111 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 io_wbs_datrd[2]
port 112 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 io_wbs_datrd[30]
port 113 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 io_wbs_datrd[31]
port 114 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_wbs_datrd[3]
port 115 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 io_wbs_datrd[4]
port 116 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 io_wbs_datrd[5]
port 117 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_wbs_datrd[6]
port 118 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 io_wbs_datrd[7]
port 119 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 io_wbs_datrd[8]
port 120 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 io_wbs_datrd[9]
port 121 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 io_wbs_datwr[0]
port 122 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 io_wbs_datwr[10]
port 123 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 io_wbs_datwr[11]
port 124 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 io_wbs_datwr[12]
port 125 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 io_wbs_datwr[13]
port 126 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 io_wbs_datwr[14]
port 127 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 io_wbs_datwr[15]
port 128 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 io_wbs_datwr[16]
port 129 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 io_wbs_datwr[17]
port 130 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 io_wbs_datwr[18]
port 131 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 io_wbs_datwr[19]
port 132 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_datwr[1]
port 133 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 io_wbs_datwr[20]
port 134 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 io_wbs_datwr[21]
port 135 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 io_wbs_datwr[22]
port 136 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 io_wbs_datwr[23]
port 137 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 io_wbs_datwr[24]
port 138 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 io_wbs_datwr[25]
port 139 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 io_wbs_datwr[26]
port 140 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 io_wbs_datwr[27]
port 141 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 io_wbs_datwr[28]
port 142 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 io_wbs_datwr[29]
port 143 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 io_wbs_datwr[2]
port 144 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 io_wbs_datwr[30]
port 145 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 io_wbs_datwr[31]
port 146 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 io_wbs_datwr[3]
port 147 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 io_wbs_datwr[4]
port 148 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 io_wbs_datwr[5]
port 149 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 io_wbs_datwr[6]
port 150 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 io_wbs_datwr[7]
port 151 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_wbs_datwr[8]
port 152 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 io_wbs_datwr[9]
port 153 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 io_wbs_rst
port 154 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_wbs_stb
port 155 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 io_wbs_we
port 156 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 157 nsew power input
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 157 nsew power input
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 157 nsew power input
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 157 nsew power input
rlabel metal4 s 127088 2128 127408 107760 6 vccd1
port 157 nsew power input
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 158 nsew ground input
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 158 nsew ground input
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 158 nsew ground input
rlabel metal4 s 111728 2128 112048 107760 6 vssd1
port 158 nsew ground input
rlabel metal4 s 142448 2128 142768 107760 6 vssd1
port 158 nsew ground input
rlabel metal2 s 11334 109200 11390 110000 6 wfg_drive_pat_dout_o[0]
port 159 nsew signal output
rlabel metal2 s 43902 109200 43958 110000 6 wfg_drive_pat_dout_o[10]
port 160 nsew signal output
rlabel metal2 s 47214 109200 47270 110000 6 wfg_drive_pat_dout_o[11]
port 161 nsew signal output
rlabel metal2 s 50434 109200 50490 110000 6 wfg_drive_pat_dout_o[12]
port 162 nsew signal output
rlabel metal2 s 53654 109200 53710 110000 6 wfg_drive_pat_dout_o[13]
port 163 nsew signal output
rlabel metal2 s 56966 109200 57022 110000 6 wfg_drive_pat_dout_o[14]
port 164 nsew signal output
rlabel metal2 s 60186 109200 60242 110000 6 wfg_drive_pat_dout_o[15]
port 165 nsew signal output
rlabel metal2 s 63498 109200 63554 110000 6 wfg_drive_pat_dout_o[16]
port 166 nsew signal output
rlabel metal2 s 66718 109200 66774 110000 6 wfg_drive_pat_dout_o[17]
port 167 nsew signal output
rlabel metal2 s 70030 109200 70086 110000 6 wfg_drive_pat_dout_o[18]
port 168 nsew signal output
rlabel metal2 s 73250 109200 73306 110000 6 wfg_drive_pat_dout_o[19]
port 169 nsew signal output
rlabel metal2 s 14554 109200 14610 110000 6 wfg_drive_pat_dout_o[1]
port 170 nsew signal output
rlabel metal2 s 76562 109200 76618 110000 6 wfg_drive_pat_dout_o[20]
port 171 nsew signal output
rlabel metal2 s 79782 109200 79838 110000 6 wfg_drive_pat_dout_o[21]
port 172 nsew signal output
rlabel metal2 s 83002 109200 83058 110000 6 wfg_drive_pat_dout_o[22]
port 173 nsew signal output
rlabel metal2 s 86314 109200 86370 110000 6 wfg_drive_pat_dout_o[23]
port 174 nsew signal output
rlabel metal2 s 89534 109200 89590 110000 6 wfg_drive_pat_dout_o[24]
port 175 nsew signal output
rlabel metal2 s 92846 109200 92902 110000 6 wfg_drive_pat_dout_o[25]
port 176 nsew signal output
rlabel metal2 s 96066 109200 96122 110000 6 wfg_drive_pat_dout_o[26]
port 177 nsew signal output
rlabel metal2 s 99378 109200 99434 110000 6 wfg_drive_pat_dout_o[27]
port 178 nsew signal output
rlabel metal2 s 102598 109200 102654 110000 6 wfg_drive_pat_dout_o[28]
port 179 nsew signal output
rlabel metal2 s 105818 109200 105874 110000 6 wfg_drive_pat_dout_o[29]
port 180 nsew signal output
rlabel metal2 s 17866 109200 17922 110000 6 wfg_drive_pat_dout_o[2]
port 181 nsew signal output
rlabel metal2 s 109130 109200 109186 110000 6 wfg_drive_pat_dout_o[30]
port 182 nsew signal output
rlabel metal2 s 112350 109200 112406 110000 6 wfg_drive_pat_dout_o[31]
port 183 nsew signal output
rlabel metal2 s 21086 109200 21142 110000 6 wfg_drive_pat_dout_o[3]
port 184 nsew signal output
rlabel metal2 s 24398 109200 24454 110000 6 wfg_drive_pat_dout_o[4]
port 185 nsew signal output
rlabel metal2 s 27618 109200 27674 110000 6 wfg_drive_pat_dout_o[5]
port 186 nsew signal output
rlabel metal2 s 30838 109200 30894 110000 6 wfg_drive_pat_dout_o[6]
port 187 nsew signal output
rlabel metal2 s 34150 109200 34206 110000 6 wfg_drive_pat_dout_o[7]
port 188 nsew signal output
rlabel metal2 s 37370 109200 37426 110000 6 wfg_drive_pat_dout_o[8]
port 189 nsew signal output
rlabel metal2 s 40682 109200 40738 110000 6 wfg_drive_pat_dout_o[9]
port 190 nsew signal output
rlabel metal2 s 1582 109200 1638 110000 6 wfg_drive_spi_cs_no
port 191 nsew signal output
rlabel metal2 s 4802 109200 4858 110000 6 wfg_drive_spi_sclk_o
port 192 nsew signal output
rlabel metal2 s 8022 109200 8078 110000 6 wfg_drive_spi_sdo_o
port 193 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 150000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36007748
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/wfg/runs/wfg/results/finishing/wfg_top.magic.gds
string GDS_START 1586680
<< end >>

