magic
tech sky130A
magscale 1 2
timestamp 1657783272
<< nwell >>
rect 1066 37253 118902 37574
rect 1066 36165 118902 36731
rect 1066 35077 118902 35643
rect 1066 33989 118902 34555
rect 1066 32901 118902 33467
rect 1066 31813 118902 32379
rect 1066 30725 118902 31291
rect 1066 29637 118902 30203
rect 1066 28549 118902 29115
rect 1066 27461 118902 28027
rect 1066 26373 118902 26939
rect 1066 25285 118902 25851
rect 1066 24197 118902 24763
rect 1066 23109 118902 23675
rect 1066 22021 118902 22587
rect 1066 20933 118902 21499
rect 1066 19845 118902 20411
rect 1066 18757 118902 19323
rect 1066 17669 118902 18235
rect 1066 16581 118902 17147
rect 1066 15493 118902 16059
rect 1066 14405 118902 14971
rect 1066 13317 118902 13883
rect 1066 12229 118902 12795
rect 1066 11141 118902 11707
rect 1066 10053 118902 10619
rect 1066 8965 118902 9531
rect 1066 7877 118902 8443
rect 1066 6789 118902 7355
rect 1066 5701 118902 6267
rect 1066 4613 118902 5179
rect 1066 3525 118902 4091
rect 1066 2437 118902 3003
<< obsli1 >>
rect 1104 2159 118864 37553
<< obsm1 >>
rect 1104 484 118864 37584
<< metal2 >>
rect 2686 0 2742 800
rect 4066 0 4122 800
rect 5446 0 5502 800
rect 6826 0 6882 800
rect 8206 0 8262 800
rect 9586 0 9642 800
rect 10966 0 11022 800
rect 12346 0 12402 800
rect 13726 0 13782 800
rect 15106 0 15162 800
rect 16486 0 16542 800
rect 17866 0 17922 800
rect 19246 0 19302 800
rect 20626 0 20682 800
rect 22006 0 22062 800
rect 23386 0 23442 800
rect 24766 0 24822 800
rect 26146 0 26202 800
rect 27526 0 27582 800
rect 28906 0 28962 800
rect 30286 0 30342 800
rect 31666 0 31722 800
rect 33046 0 33102 800
rect 34426 0 34482 800
rect 35806 0 35862 800
rect 37186 0 37242 800
rect 38566 0 38622 800
rect 39946 0 40002 800
rect 41326 0 41382 800
rect 42706 0 42762 800
rect 44086 0 44142 800
rect 45466 0 45522 800
rect 46846 0 46902 800
rect 48226 0 48282 800
rect 49606 0 49662 800
rect 50986 0 51042 800
rect 52366 0 52422 800
rect 53746 0 53802 800
rect 55126 0 55182 800
rect 56506 0 56562 800
rect 57886 0 57942 800
rect 59266 0 59322 800
rect 60646 0 60702 800
rect 62026 0 62082 800
rect 63406 0 63462 800
rect 64786 0 64842 800
rect 66166 0 66222 800
rect 67546 0 67602 800
rect 68926 0 68982 800
rect 70306 0 70362 800
rect 71686 0 71742 800
rect 73066 0 73122 800
rect 74446 0 74502 800
rect 75826 0 75882 800
rect 77206 0 77262 800
rect 78586 0 78642 800
rect 79966 0 80022 800
rect 81346 0 81402 800
rect 82726 0 82782 800
rect 84106 0 84162 800
rect 85486 0 85542 800
rect 86866 0 86922 800
rect 88246 0 88302 800
rect 89626 0 89682 800
rect 91006 0 91062 800
rect 92386 0 92442 800
rect 93766 0 93822 800
rect 95146 0 95202 800
rect 96526 0 96582 800
rect 97906 0 97962 800
rect 99286 0 99342 800
rect 100666 0 100722 800
rect 102046 0 102102 800
rect 103426 0 103482 800
rect 104806 0 104862 800
rect 106186 0 106242 800
rect 107566 0 107622 800
rect 108946 0 109002 800
rect 110326 0 110382 800
rect 111706 0 111762 800
rect 113086 0 113142 800
rect 114466 0 114522 800
rect 115846 0 115902 800
rect 117226 0 117282 800
<< obsm2 >>
rect 2688 856 118202 37573
rect 2798 478 4010 856
rect 4178 478 5390 856
rect 5558 478 6770 856
rect 6938 478 8150 856
rect 8318 478 9530 856
rect 9698 478 10910 856
rect 11078 478 12290 856
rect 12458 478 13670 856
rect 13838 478 15050 856
rect 15218 478 16430 856
rect 16598 478 17810 856
rect 17978 478 19190 856
rect 19358 478 20570 856
rect 20738 478 21950 856
rect 22118 478 23330 856
rect 23498 478 24710 856
rect 24878 478 26090 856
rect 26258 478 27470 856
rect 27638 478 28850 856
rect 29018 478 30230 856
rect 30398 478 31610 856
rect 31778 478 32990 856
rect 33158 478 34370 856
rect 34538 478 35750 856
rect 35918 478 37130 856
rect 37298 478 38510 856
rect 38678 478 39890 856
rect 40058 478 41270 856
rect 41438 478 42650 856
rect 42818 478 44030 856
rect 44198 478 45410 856
rect 45578 478 46790 856
rect 46958 478 48170 856
rect 48338 478 49550 856
rect 49718 478 50930 856
rect 51098 478 52310 856
rect 52478 478 53690 856
rect 53858 478 55070 856
rect 55238 478 56450 856
rect 56618 478 57830 856
rect 57998 478 59210 856
rect 59378 478 60590 856
rect 60758 478 61970 856
rect 62138 478 63350 856
rect 63518 478 64730 856
rect 64898 478 66110 856
rect 66278 478 67490 856
rect 67658 478 68870 856
rect 69038 478 70250 856
rect 70418 478 71630 856
rect 71798 478 73010 856
rect 73178 478 74390 856
rect 74558 478 75770 856
rect 75938 478 77150 856
rect 77318 478 78530 856
rect 78698 478 79910 856
rect 80078 478 81290 856
rect 81458 478 82670 856
rect 82838 478 84050 856
rect 84218 478 85430 856
rect 85598 478 86810 856
rect 86978 478 88190 856
rect 88358 478 89570 856
rect 89738 478 90950 856
rect 91118 478 92330 856
rect 92498 478 93710 856
rect 93878 478 95090 856
rect 95258 478 96470 856
rect 96638 478 97850 856
rect 98018 478 99230 856
rect 99398 478 100610 856
rect 100778 478 101990 856
rect 102158 478 103370 856
rect 103538 478 104750 856
rect 104918 478 106130 856
rect 106298 478 107510 856
rect 107678 478 108890 856
rect 109058 478 110270 856
rect 110438 478 111650 856
rect 111818 478 113030 856
rect 113198 478 114410 856
rect 114578 478 115790 856
rect 115958 478 117170 856
rect 117338 478 118202 856
<< metal3 >>
rect 119200 37000 120000 37120
rect 119200 36184 120000 36304
rect 119200 35368 120000 35488
rect 119200 34552 120000 34672
rect 119200 33736 120000 33856
rect 119200 32920 120000 33040
rect 119200 32104 120000 32224
rect 119200 31288 120000 31408
rect 119200 30472 120000 30592
rect 119200 29656 120000 29776
rect 119200 28840 120000 28960
rect 119200 28024 120000 28144
rect 119200 27208 120000 27328
rect 119200 26392 120000 26512
rect 119200 25576 120000 25696
rect 119200 24760 120000 24880
rect 119200 23944 120000 24064
rect 119200 23128 120000 23248
rect 119200 22312 120000 22432
rect 119200 21496 120000 21616
rect 119200 20680 120000 20800
rect 119200 19864 120000 19984
rect 119200 19048 120000 19168
rect 119200 18232 120000 18352
rect 119200 17416 120000 17536
rect 119200 16600 120000 16720
rect 119200 15784 120000 15904
rect 119200 14968 120000 15088
rect 119200 14152 120000 14272
rect 119200 13336 120000 13456
rect 119200 12520 120000 12640
rect 119200 11704 120000 11824
rect 119200 10888 120000 11008
rect 119200 10072 120000 10192
rect 119200 9256 120000 9376
rect 119200 8440 120000 8560
rect 119200 7624 120000 7744
rect 119200 6808 120000 6928
rect 119200 5992 120000 6112
rect 119200 5176 120000 5296
rect 119200 4360 120000 4480
rect 119200 3544 120000 3664
rect 119200 2728 120000 2848
<< obsm3 >>
rect 4210 37200 119200 37569
rect 4210 36920 119120 37200
rect 4210 36384 119200 36920
rect 4210 36104 119120 36384
rect 4210 35568 119200 36104
rect 4210 35288 119120 35568
rect 4210 34752 119200 35288
rect 4210 34472 119120 34752
rect 4210 33936 119200 34472
rect 4210 33656 119120 33936
rect 4210 33120 119200 33656
rect 4210 32840 119120 33120
rect 4210 32304 119200 32840
rect 4210 32024 119120 32304
rect 4210 31488 119200 32024
rect 4210 31208 119120 31488
rect 4210 30672 119200 31208
rect 4210 30392 119120 30672
rect 4210 29856 119200 30392
rect 4210 29576 119120 29856
rect 4210 29040 119200 29576
rect 4210 28760 119120 29040
rect 4210 28224 119200 28760
rect 4210 27944 119120 28224
rect 4210 27408 119200 27944
rect 4210 27128 119120 27408
rect 4210 26592 119200 27128
rect 4210 26312 119120 26592
rect 4210 25776 119200 26312
rect 4210 25496 119120 25776
rect 4210 24960 119200 25496
rect 4210 24680 119120 24960
rect 4210 24144 119200 24680
rect 4210 23864 119120 24144
rect 4210 23328 119200 23864
rect 4210 23048 119120 23328
rect 4210 22512 119200 23048
rect 4210 22232 119120 22512
rect 4210 21696 119200 22232
rect 4210 21416 119120 21696
rect 4210 20880 119200 21416
rect 4210 20600 119120 20880
rect 4210 20064 119200 20600
rect 4210 19784 119120 20064
rect 4210 19248 119200 19784
rect 4210 18968 119120 19248
rect 4210 18432 119200 18968
rect 4210 18152 119120 18432
rect 4210 17616 119200 18152
rect 4210 17336 119120 17616
rect 4210 16800 119200 17336
rect 4210 16520 119120 16800
rect 4210 15984 119200 16520
rect 4210 15704 119120 15984
rect 4210 15168 119200 15704
rect 4210 14888 119120 15168
rect 4210 14352 119200 14888
rect 4210 14072 119120 14352
rect 4210 13536 119200 14072
rect 4210 13256 119120 13536
rect 4210 12720 119200 13256
rect 4210 12440 119120 12720
rect 4210 11904 119200 12440
rect 4210 11624 119120 11904
rect 4210 11088 119200 11624
rect 4210 10808 119120 11088
rect 4210 10272 119200 10808
rect 4210 9992 119120 10272
rect 4210 9456 119200 9992
rect 4210 9176 119120 9456
rect 4210 8640 119200 9176
rect 4210 8360 119120 8640
rect 4210 7824 119200 8360
rect 4210 7544 119120 7824
rect 4210 7008 119200 7544
rect 4210 6728 119120 7008
rect 4210 6192 119200 6728
rect 4210 5912 119120 6192
rect 4210 5376 119200 5912
rect 4210 5096 119120 5376
rect 4210 4560 119200 5096
rect 4210 4280 119120 4560
rect 4210 3744 119200 4280
rect 4210 3464 119120 3744
rect 4210 2928 119200 3464
rect 4210 2648 119120 2928
rect 4210 1123 119200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
rect 111728 2128 112048 37584
<< labels >>
rlabel metal3 s 119200 3544 120000 3664 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 119200 4360 120000 4480 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 119200 5176 120000 5296 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 119200 5992 120000 6112 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 119200 7624 120000 7744 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 119200 8440 120000 8560 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 119200 9256 120000 9376 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 119200 10072 120000 10192 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 119200 10888 120000 11008 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 119200 2728 120000 2848 6 csb
port 29 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 119200 11704 120000 11824 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 119200 19864 120000 19984 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 119200 20680 120000 20800 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 119200 21496 120000 21616 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 119200 22312 120000 22432 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 119200 23128 120000 23248 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 119200 23944 120000 24064 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 119200 24760 120000 24880 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 119200 25576 120000 25696 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 119200 26392 120000 26512 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 119200 27208 120000 27328 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 119200 12520 120000 12640 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 119200 28024 120000 28144 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 119200 28840 120000 28960 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 119200 29656 120000 29776 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 119200 30472 120000 30592 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 119200 31288 120000 31408 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 119200 32104 120000 32224 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 119200 32920 120000 33040 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 119200 33736 120000 33856 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 119200 34552 120000 34672 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 119200 35368 120000 35488 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 119200 13336 120000 13456 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 119200 36184 120000 36304 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 119200 37000 120000 37120 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 119200 14152 120000 14272 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 119200 14968 120000 15088 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 119200 15784 120000 15904 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 119200 16600 120000 16720 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 119200 17416 120000 17536 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 119200 18232 120000 18352 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 119200 19048 120000 19168 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 129 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1616618
string GDS_FILE /home/leo/Dokumente/caravel_workspace_mpw7/caravel_wfg/openlane/merge_memory/runs/22_07_14_09_20/results/signoff/merge_memory.magic.gds
string GDS_START 51508
<< end >>

